VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO AssuraMatchStatus STRING ;
  MACRO connectivityLastUpdated INTEGER ;
  MACRO _mspsExtractedMode STRING ;
  MACRO _mspsExtractionCreatedBy STRING ;
  MACRO extractionCreatedBy STRING ;
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_WIDTH STRING ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.01 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER NWEL
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
  PROPERTY LEF58_SPACING "SPACING 2.2 ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.9 ;" ;
END NWEL

LAYER DIFF
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE DIFFUSION ;" ;
  PROPERTY LEF58_SPACING "SPACING 0.28 ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.24 ;" ;
END DIFF

LAYER PPLUS
  TYPE IMPLANT ;
  WIDTH 0.4 ;
  SPACING 0.4 ;
  AREA 0.2916 ;
END PPLUS

LAYER NPLUS
  TYPE IMPLANT ;
  WIDTH 0.4 ;
  SPACING 0.4 ;
  AREA 0.2916 ;
END NPLUS

LAYER PO1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.18 ;
  AREA 0.198 ;
  SPACING 0.34 ;
  RESISTANCE RPERSQ 8 ;
  PROPERTY LEF58_TYPE "TYPE POLYROUTING ;" ;
END PO1

LAYER CONT
  TYPE CUT ;
  SPACING 0.26 ;
  WIDTH 0.24 ;
  ENCLOSURE BELOW 0.1 0.1 ;
  ENCLOSURE ABOVE 0 0.08 ;
END CONT

LAYER ME1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.48 0.48 ;
  WIDTH 0.24 ;
  OFFSET 0.24 0.24 ;
  AREA 0.1764 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 9.999 
    WIDTH 0 0.24 0.28 
    WIDTH 9.999 0.28 0.28 ;
  RESISTANCE RPERSQ 0.077 ;
  MINIMUMDENSITY 25 ;
  DENSITYCHECKWINDOW 1000 1000 ;
  DENSITYCHECKSTEP 500 ;
END ME1

LAYER VI1
  TYPE CUT ;
  SPACING 0.28 ;
  WIDTH 0.28 ;
  ENCLOSURE BELOW 0.2 0.08 WIDTH 10 ;
  ENCLOSURE BELOW 0 0.08 ;
  ENCLOSURE ABOVE 0 0.08 ;
END VI1

LAYER ME2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.56 0.56 ;
  WIDTH 0.28 ;
  OFFSET 0.28 0.28 ;
  AREA 0.1936 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 9.999 
    WIDTH 0 0.28 0.32 
    WIDTH 9.999 0.32 0.32 ;
  RESISTANCE RPERSQ 0.062 ;
  MINIMUMDENSITY 25 ;
  DENSITYCHECKWINDOW 1000 1000 ;
  DENSITYCHECKSTEP 500 ;
END ME2

LAYER VI2
  TYPE CUT ;
  SPACING 0.28 ;
  WIDTH 0.28 ;
  ENCLOSURE BELOW 0.2 0.08 WIDTH 10 ;
  ENCLOSURE BELOW 0 0.08 ;
  ENCLOSURE ABOVE 0 0.08 ;
END VI2

LAYER ME3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.56 0.56 ;
  WIDTH 0.28 ;
  OFFSET 0.28 0.28 ;
  AREA 0.1936 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 9.999 
    WIDTH 0 0.28 0.32 
    WIDTH 9.999 0.32 0.32 ;
  RESISTANCE RPERSQ 0.062 ;
  MINIMUMDENSITY 25 ;
  DENSITYCHECKWINDOW 1000 1000 ;
  DENSITYCHECKSTEP 500 ;
END ME3

LAYER VI3
  TYPE CUT ;
  SPACING 0.28 ;
  WIDTH 0.28 ;
  ENCLOSURE BELOW 0.2 0.08 WIDTH 10 ;
  ENCLOSURE BELOW 0 0.08 ;
  ENCLOSURE ABOVE 0 0.08 ;
END VI3

LAYER ME4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.56 0.56 ;
  WIDTH 0.28 ;
  OFFSET 0.28 0.28 ;
  AREA 0.1936 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 9.999 
    WIDTH 0 0.28 0.32 
    WIDTH 9.999 0.32 0.32 ;
  RESISTANCE RPERSQ 0.062 ;
  MINIMUMDENSITY 25 ;
  DENSITYCHECKWINDOW 1000 1000 ;
  DENSITYCHECKSTEP 500 ;
END ME4

LAYER VI4
  TYPE CUT ;
  SPACING 0.28 ;
  WIDTH 0.28 ;
  ENCLOSURE BELOW 0.2 0.08 WIDTH 10 ;
  ENCLOSURE BELOW 0 0.08 ;
  ENCLOSURE ABOVE 0 0.08 ;
END VI4

LAYER ME5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.56 0.56 ;
  WIDTH 0.28 ;
  OFFSET 0.28 0.28 ;
  AREA 0.1936 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 9.999 
    WIDTH 0 0.28 0.32 
    WIDTH 9.999 0.32 0.32 ;
  RESISTANCE RPERSQ 0.062 ;
  MINIMUMDENSITY 25 ;
  DENSITYCHECKWINDOW 1000 1000 ;
  DENSITYCHECKSTEP 500 ;
END ME5

LAYER VI5
  TYPE CUT ;
  SPACING 0.28 ;
  WIDTH 0.28 ;
  ENCLOSURE BELOW 0.2 0.08 WIDTH 10 ;
  ENCLOSURE BELOW 0 0.08 ;
  ENCLOSURE ABOVE 0.4 0.4 ;
END VI5

LAYER ME6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 2.2 2.2 ;
  WIDTH 1.2 ;
  OFFSET 1.1 1.1 ;
  AREA 9 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 9.999 
    WIDTH 0 1 1.5 
    WIDTH 9.999 1.5 1.5 ;
  RESISTANCE RPERSQ 0.02 ;
  MINIMUMDENSITY 25 ;
  DENSITYCHECKWINDOW 1000 1000 ;
  DENSITYCHECKSTEP 500 ;
END ME6

VIARULE M5_M6 GENERATE DEFAULT
  LAYER ME5 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER ME6 ;
    ENCLOSURE 0.4 0.4 ;
  LAYER VI5 ;
    RECT -0.14 -0.14 0.14 0.14 ;
    SPACING 0.56 BY 0.56 ;
END M5_M6

VIARULE M4_M5 GENERATE DEFAULT
  LAYER ME4 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER ME5 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER VI4 ;
    RECT -0.14 -0.14 0.14 0.14 ;
    SPACING 0.56 BY 0.56 ;
END M4_M5

VIARULE M3_M4 GENERATE DEFAULT
  LAYER ME3 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER ME4 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER VI3 ;
    RECT -0.14 -0.14 0.14 0.14 ;
    SPACING 0.56 BY 0.56 ;
END M3_M4

VIARULE M2_M3 GENERATE DEFAULT
  LAYER ME2 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER ME3 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER VI2 ;
    RECT -0.14 -0.14 0.14 0.14 ;
    SPACING 0.56 BY 0.56 ;
END M2_M3

VIARULE M1_M2 GENERATE DEFAULT
  LAYER ME1 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER ME2 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER VI1 ;
    RECT -0.14 -0.14 0.14 0.14 ;
    SPACING 0.56 BY 0.56 ;
END M1_M2

VIARULE M1_PDIFF GENERATE
  LAYER DIFF ;
    ENCLOSURE 0.1 0.1 ;
  LAYER ME1 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER CONT ;
    RECT -0.12 -0.12 0.12 0.12 ;
    SPACING 0.5 BY 0.5 ;
END M1_PDIFF

VIARULE M1_NWEL GENERATE
  LAYER DIFF ;
    ENCLOSURE 0.1 0.1 ;
  LAYER ME1 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER CONT ;
    RECT -0.12 -0.12 0.12 0.12 ;
    SPACING 0.5 BY 0.5 ;
END M1_NWEL

VIARULE M1_NDIFF GENERATE
  LAYER DIFF ;
    ENCLOSURE 0.1 0.1 ;
  LAYER ME1 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER CONT ;
    RECT -0.12 -0.12 0.12 0.12 ;
    SPACING 0.5 BY 0.5 ;
END M1_NDIFF

VIARULE M1_POLY GENERATE DEFAULT
  LAYER PO1 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER ME1 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER CONT ;
    RECT -0.12 -0.12 0.12 0.12 ;
    SPACING 0.5 BY 0.5 ;
END M1_POLY

MACRO AND2X1
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 8.44 0.24 8.68 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 2.73 0.24 2.97 ;
    END
  END b
  PIN y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 11.17 5.59 11.41 5.83 ;
    END
  END y
  PIN vdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 11.17 11.412 11.41 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 0 11.412 0.24 ;
    END
  END gnd
  PROPERTY AssuraMatchStatus "fully_matched" ;
  PROPERTY connectivityLastUpdated 560 ;
  PROPERTY _mspsExtractedMode "analog" ;
  PROPERTY _mspsExtractionCreatedBy "Assura" ;
  PROPERTY extractionCreatedBy "Assura" ;
END AND2X1

MACRO INVX1
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 3.16 0.24 3.4 ;
    END
  END a
  PIN vdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 6.32 6.56 6.56 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 0 6.56 0.24 ;
    END
  END gnd
  PIN y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 6.32 3.16 6.56 3.4 ;
    END
  END y
  PROPERTY AssuraMatchStatus "fully_matched" ;
  PROPERTY connectivityLastUpdated 287 ;
  PROPERTY _mspsExtractedMode "analog" ;
  PROPERTY _mspsExtractionCreatedBy "Assura" ;
  PROPERTY extractionCreatedBy "Assura" ;
END INVX1

MACRO NAND2X1
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 6.92 0.24 7.16 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 2.23 0.24 2.47 ;
    END
  END b
  PIN y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 9.14 4.57 9.38 4.81 ;
    END
  END y
  PIN vdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 9.14 9.385 9.38 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 0 9.385 0.24 ;
    END
  END gnd
  PROPERTY AssuraMatchStatus "fully_matched" ;
  PROPERTY connectivityLastUpdated 676 ;
  PROPERTY _mspsExtractedMode "analog" ;
  PROPERTY _mspsExtractionCreatedBy "Assura" ;
  PROPERTY extractionCreatedBy "Assura" ;
END NAND2X1

MACRO NOR2X1
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 7.7 0.24 7.94 ;
    END
  END a
  PIN y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 10.18 5.09 10.42 5.33 ;
    END
  END y
  PIN gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 0 10.427 0.24 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 10.18 10.427 10.42 ;
    END
  END vdd
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 2.49 0.24 2.73 ;
    END
  END b
  PROPERTY AssuraMatchStatus "fully_matched" ;
  PROPERTY connectivityLastUpdated 686 ;
  PROPERTY _mspsExtractedMode "analog" ;
  PROPERTY _mspsExtractionCreatedBy "Assura" ;
  PROPERTY extractionCreatedBy "Assura" ;
END NOR2X1

MACRO OR2X1
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 9.09 0.24 9.33 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 2.95 0.24 3.19 ;
    END
  END b
  PIN y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 12.04 6.02 12.28 6.26 ;
    END
  END y
  PIN vdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 12.04 12.283 12.28 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 0 0 12.283 0.24 ;
    END
  END gnd
  PROPERTY AssuraMatchStatus "fully_matched" ;
  PROPERTY connectivityLastUpdated 1052 ;
  PROPERTY _mspsExtractedMode "analog" ;
  PROPERTY _mspsExtractionCreatedBy "Assura" ;
  PROPERTY extractionCreatedBy "Assura" ;
END OR2X1

END LIBRARY
