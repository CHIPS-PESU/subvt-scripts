*
*
*
*                       LINUX           Tue May 18 23:28:51 2021
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus - (64-bit)
*  Version        : 20.1.1-s233
*  Build Date     : Wed Mar 25 13:13:47 PDT 2020
*
*  HSPICE LIBRARY
*
*
*

*
.SUBCKT XOR2X1 vdd gnd a b y
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
M9	vdd#3	a#13	gnd#3	gnd#11	n_18_mm	L=1.8e-07
+ W=2.4e-07	effW=2.4e-07
M10	net12#3	b#7	gnd#14	gnd#11	n_18_mm
+ L=1.8e-07	W=2.4e-07
+ effW=2.4e-07
M4	y#8	a#10	net29#2	gnd#11	n_18_mm
+ L=1.8e-07	W=4.8e-07
+ effW=4.8e-07
M6	net29	b#5	gnd#13	gnd#11	n_18_mm
+ L=1.8e-07	W=4.8e-07
+ effW=4.8e-07
M5	y#5	vdd#13	net28	gnd#11	n_18_mm
+ L=1.8e-07	W=4.8e-07
+ effW=4.8e-07
M7	net28#3	net12#16	gnd#7	gnd#11	n_18_mm
+ L=1.8e-07	W=4.8e-07
+ effW=4.8e-07
M8	vdd#49	a#14	vdd#1	vdd#34	p_18_mm
+ L=1.8e-07	W=3.18e-06
+ effW=3.18e-06
M11	net12#4	b#8	vdd#50	vdd#38	p_18_mm
+ L=1.8e-07	W=3.18e-06
+ effW=3.18e-06
M0	net31#3	a#8	vdd#48	vdd#41	p_18_mm
+ L=1.8e-07	W=3.18e-06
+ effW=3.18e-06
M2	y#1	net12#12	net31#6	vdd#45	p_18_mm
+ L=1.8e-07	W=3.18e-06
+ effW=3.18e-06
M0@1	net31#3	a#11	vdd#47	vdd#41	p_18_mm
+ L=1.8e-07	W=3.18e-06
+ effW=3.18e-06
M2@1	y#1	net12#9	net31	vdd#45	p_18_mm
+ L=1.8e-07	W=3.18e-06
+ effW=3.18e-06
MavD28_7_unmatched	vdd#9	vdd#28	vdd#40	vdd#41
+ p_18_mm	L=1.8e-07	W=3.18e-06	effW=3.18e-06
MavD28_8_unmatched	y#10	b#10	vdd#17	vdd#45	p_18_mm
+ L=1.8e-07	W=3.18e-06
+ effW=3.18e-06
MavD28_9_unmatched	vdd#18	vdd#24	vdd#9	vdd#41
+ p_18_mm	L=1.8237e-07	W=3.38e-06	effW=3.38e-06
MavD28_10_unmatched	vdd#15	avC10	y#10	vdd#45	p_18_mm
+ L=1.8157e-07	W=3.31e-06
+ effW=3.31e-06
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rh1	a#8	a#6	  105.0147	$PLY_C
Rh2	a#10	a#9	   24.9369	$PLY_C
Rh3	a#11	a#5	  211.9010	$PLY_C
Rh4	a#5	a#3	   82.8930	$PLY_C
Rh5	a#3	a#12	    2.9102	$PLY_C
Rh6	a#12	a#1	  194.1718	$PLY_C
Rh7	a#3	a#13	   27.8774	$PLY_C
Rh8	a#12	a#2	   41.6306	$PLY_C
Rh9	a#2	a#14	   84.9368	$PLY_C
Rh10	net12#9	net12#10	  108.9094	$PLY_C
Rh11	net12#10	net12#11	   37.0830	$PLY_C
Rh12	net12#11	net12#8	    5.2372	$PLY_C
Rh13	net12#10	net12#12	   77.6199	$PLY_C
Rh14	net12#11	net12#13	   40.8895	$PLY_C
Rh15	b#5	b#4	   23.6888	$PLY_C
Rh16	b#4	b#3	  139.0704	$PLY_C
Rh17	b#3	b#2	   28.7110	$PLY_C
Rh18	b#2	b#1	  205.3490	$PLY_C
Rh19	b#4	b#6	  234.8601	$PLY_C
Rh20	b#3	b#7	   27.4666	$PLY_C
Rh21	b#2	b#8	   83.6376	$PLY_C
Rh22	b#10	b#9	  105.0147	$PLY_C
Rh23	vdd#13	vdd#14	   36.9369	$PLY_C
Rh24	net12#16	net12#15	   23.6888	$PLY_C
Rh25	net12#15	net12#14	  181.2188	$PLY_C
Rh26	vdd#24	vdd#25	   66.3887	$PLY_C
Rh27	vdd#25	vdd#20	    2.3662	$PLY_C
Rh28	vdd#20	vdd#26	   19.6286	$PLY_C
Rh29	vdd#26	vdd#6	   44.9074	$PLY_C
Rh30	vdd#26	vdd#28	   71.9261	$PLY_C
Rh31	vdd#8	vdd#25	   12.0000	$PLY_C
Rg1	b	b#1	   12.2018	$ME1_C
Rg2	a#1	a	   12.9240	$ME1_C
Rg3	gnd#1	gnd#2	4.596e-03	$ME1_C
Rg4	gnd#4	gnd#5	4.596e-03	$ME1_C
Rg5	gnd#1	gnd#5	9.704e-02	$ME1_C
Rg6	gnd#3	gnd#4	   15.0000	$ME1_C
Rg7	net12#3	net12#5	   16.1506	$ME1_C
Rg8	net12#5	net12#2	    0.5424	$ME1_C
Rg9	net12#4	net12#5	    2.5000	$ME1_C
Rg10	vdd#1	vdd#2	    2.6464	$ME1_C
Rg11	vdd#2	vdd#3	   16.0609	$ME1_C
Rg12	vdd#2	vdd#4	    6.9956	$ME1_C
Rg13	net12#8	net12#7	   12.2027	$ME1_C
Rg14	a#4	a#5	   12.3353	$ME1_C
Rg15	a#4	a#6	   12.1300	$ME1_C
Rg16	a#9	a#7	   12.4031	$ME1_C
Rg17	y#1	y#2	    9.1766	$ME1_C
Rg18	net29	net29#3	   15.8650	$ME1_C
Rg19	net29#3	net29#2	   15.0214	$ME1_C
Rg20	net29#2	net29#3	   15.0000	$ME1_C
Rg21	net31	net31#2	    3.5089	$ME1_C
Rg22	net31#2	net31#4	    0.2059	$ME1_C
Rg23	net31#4	net31#5	1.941e-03	$ME1_C
Rg24	net31#2	net31#6	    3.4062	$ME1_C
Rg25	net31#5	net31#3	    3.2892	$ME1_C
Rg26	net31#3	net31#4	   15.0000	$ME1_C
Rg27	net31#3	net31#5	   15.0000	$ME1_C
Rg28	b#9	b#6	   12.3016	$ME1_C
Rg29	net12#14	net12#13	   13.1100	$ME1_C
Rg30	y#4	y#6	1.060e-02	$ME1_C
Rg31	y#6	y#7	    0.6530	$ME1_C
Rg32	y#7	y#8	   15.2609	$ME1_C
Rg33	y#7	y#3	    0.3274	$ME1_C
Rg34	y#5	y#6	   15.0000	$ME1_C
Rg35	vdd#8	vdd#10	1.261e-02	$ME1_C
Rg36	vdd#10	vdd#11	8.733e-03	$ME1_C
Rg37	vdd#11	vdd#12	    0.2746	$ME1_C
Rg38	vdd#12	vdd#9	    3.0011	$ME1_C
Rg39	vdd#9	vdd#10	   15.0000	$ME1_C
Rg40	vdd#9	vdd#11	   15.0000	$ME1_C
Rg41	y#9	y#10	    9.2368	$ME1_C
Rg42	net28	net28#2	   15.0214	$ME1_C
Rg43	net28#2	net28#3	   15.8497	$ME1_C
Rg44	net28	net28#2	   15.0000	$ME1_C
Rg45	vdd#15	vdd#16	    3.1748	$ME1_C
Rg46	vdd#16	vdd#17	    3.2647	$ME1_C
Rg47	vdd#19	vdd#20	    6.1380	$ME1_C
Rg48	vdd#19	vdd#21	    6.8824	$ME1_C
Rg49	vdd#18	vdd#19	   15.0000	$ME1_C
Rg50	vdd#22	vdd#23	    7.3614	$ME1_C
Rg51	vdd#23	vdd#7	    0.1748	$ME1_C
Rg52	vdd#7	vdd#5	    0.8802	$ME1_C
Rg53	vdd#23	vdd#14	    0.5618	$ME1_C
Rg54	y	y#12	    1.2261	$ME1_C
Rg55	gnd#7	gnd#8	   15.3504	$ME1_C
Rg56	gnd#8	gnd	    1.2267	$ME1_C
Rg57	gnd	gnd#9	    0.1950	$ME1_C
Rg58	gnd#9	gnd#10	    0.8442	$ME1_C
Rg59	gnd#10	gnd#6	    0.5650	$ME1_C
Rg60	gnd#8	gnd#12	    1.6487	$ME1_C
Rg61	gnd#12	gnd#11	   15.0000	$ME1_C
Rg62	gnd#9	gnd#13	   15.3504	$ME1_C
Rg63	gnd#10	gnd#14	   15.3320	$ME1_C
Rg64	gnd#11	gnd#12	   15.0000	$ME1_C
Rg65	vdd#18	vdd#29	    3.7091	$ME1_C
Rg66	vdd#29	vdd#30	    0.3493	$ME1_C
Rg67	vdd#30	vdd#31	    0.3493	$ME1_C
Rg68	vdd#31	vdd	    0.1424	$ME1_C
Rg69	vdd	vdd#32	    0.3105	$ME1_C
Rg70	vdd#32	vdd#33	    0.9822	$ME1_C
Rg71	vdd#33	vdd#35	    3.2236	$ME1_C
Rg73	vdd#35	vdd#37	    2.1307	$ME1_C
Rg74	vdd#37	vdd#39	    0.3419	$ME1_C
Rg75	vdd#39	vdd#38	   15.0000	$ME1_C
Rg76	vdd#29	vdd#40	    3.2686	$ME1_C
Rg77	vdd#30	vdd#42	    0.6903	$ME1_C
Rg79	vdd#42	vdd#44	    1.0238	$ME1_C
Rg80	vdd#44	vdd#46	    0.5490	$ME1_C
Rg81	vdd#46	vdd#45	   15.0000	$ME1_C
Rg82	vdd#31	vdd#47	    3.2686	$ME1_C
Rg83	vdd#32	vdd#48	    3.2686	$ME1_C
Rg84	vdd#33	vdd#49	    3.2686	$ME1_C
Rg85	vdd#37	vdd#50	    3.3630	$ME1_C
Rg86	vdd#44	vdd#6	9.931e-02	$ME1_C
Rg88	vdd#34	vdd#35	   15.0000	$ME1_C
Rg89	vdd#34	vdd#35	   15.0000	$ME1_C
Rg90	vdd#38	vdd#39	   15.0000	$ME1_C
Rg91	vdd#41	vdd#42	   15.0000	$ME1_C
Rg92	vdd#41	vdd#42	   15.0000	$ME1_C
Rg93	vdd#45	vdd#46	   15.0000	$ME1_C
Rf1	net12	net12#2	   13.1307	$ME2_C
Rf2	gnd#2	gnd#6	   14.4116	$ME2_C
Rf3	net12#6	net12#7	   13.0974	$ME2_C
Rf4	a#4	a#7	   14.3687	$ME2_C
Rf5	vdd#5	vdd#4	    8.0476	$ME2_C
Rf6	y#3	y#2	    7.0931	$ME2_C
Rf7	vdd#6	vdd#7	   14.2270	$ME2_C
Rf8	vdd#12	vdd#16	    8.4489	$ME2_C
Rf9	y#9	y#11	    0.1589	$ME2_C
Rf10	y#11	y#4	    7.4590	$ME2_C
Rf11	y#11	y#12	    6.7560	$ME2_C
Rf12	vdd#21	vdd#22	    1.2270	$ME2_C
Re1	net12#6	net12	    0.6445	$ME3_C
*
*       CAPACITOR CARDS
*
*
C1	y#9	vdd#15	2.22329e-16
C2	net31	y#1	8.1857e-18
C3	net12#8	gnd#11	5.47628e-17
C4	y#11	net31	3.43906e-18
C5	b#2	vdd#38	6.92811e-17
C6	net12#7	net31#6	7.14538e-18
C7	a#8	net31#3	2.12414e-16
C8	a#5	vdd#45	4.8705e-17
C9	vdd#47	gnd#11	1.91086e-17
C10	gnd#5	vdd#3	2.67717e-17
C11	net12#3	b#3	3.50535e-17
C12	y#4	vdd#22	1.57449e-17
C13	vdd#13	gnd#11	3.0701e-17
C14	net12#6	vdd#50	3.83528e-17
C15	a#4	gnd#11	4.35611e-17
C16	vdd#48	a#8	2.1897e-16
C17	vdd#4	net31#2	8.84092e-17
C18	gnd#2	net12#7	1.21283e-17
C19	gnd#6	b#3	1.83206e-17
C20	vdd	gnd#11	3.30824e-17
C21	b#2	gnd#11	2.0119e-16
C22	net31#3	vdd	9.25773e-18
C23	net31	b#6	1.91661e-17
C24	a#3	vdd#3	2.63866e-17
C25	net12#8	vdd#45	2.02477e-17
C26	y#3	vdd#23	7.68538e-18
C27	vdd#5	net29#2	4.77921e-18
C28	a#6	net31#2	1.31765e-17
C29	net29	y#8	1.53807e-17
C30	vdd#13	net28	6.99119e-17
C31	net12#16	gnd#11	3.90758e-17
C32	net12#6	vdd#5	6.53336e-18
C33	a#7	gnd#11	6.79567e-17
C34	net12#12	y#1	1.57199e-16
C35	y#5	vdd#13	4.8704e-17
C36	vdd#50	net12#7	3.63333e-17
C37	b#3	gnd#11	2.4159e-16
C38	vdd#16	y#9	1.28746e-16
C39	net31#6	net12#12	1.79789e-16
C40	a#2	vdd#34	3.81285e-17
C41	a#10	gnd#11	3.34557e-17
C42	gnd#14	vdd#50	1.80609e-17
C43	vdd#48	net31#3	2.942e-16
C44	vdd#4	gnd#11	7.60499e-17
C45	net29#2	net12#14	1.54072e-18
C46	net29#2	y#8	4.97195e-17
C47	net12#16	gnd#7	5.88498e-17
C48	net12#6	a#7	5.40418e-17
C49	a	gnd#11	1.33525e-16
C50	net31#2	a#5	1.12006e-16
C51	y#4	net12#15	1.23394e-17
C52	a#2	gnd#11	5.99394e-17
C53	vdd#17	y#9	2.59343e-16
C54	gnd#2	vdd#50	3.26226e-17
C55	net28#3	net12#16	4.83155e-17
C56	b#5	gnd#11	3.91011e-17
C57	net12#6	vdd#4	8.5265e-18
C58	net31#2	a#11	1.92718e-17
C59	net31	vdd#45	1.85634e-17
C60	net28	vdd#23	9.75635e-18
C61	net12#7	gnd#11	7.4675e-17
C62	gnd#2	net12#2	1.4712e-16
C63	a#14	vdd#1	1.87341e-16
C64	vdd#2	gnd#11	3.00799e-17
C65	y#4	vdd#14	1.44984e-16
C66	b	gnd#11	7.17311e-17
C67	net29#2	a#7	1.33175e-17
C68	vdd#48	gnd#11	3.12354e-17
C69	a	vdd#34	3.06844e-17
C70	vdd#49	a#14	1.94683e-16
C71	vdd#37	a#2	2.32806e-17
C72	vdd#3	a#4	2.60076e-17
C73	a#13	gnd#11	4.73446e-17
C74	gnd#6	vdd#50	1.25005e-17
C75	y	gnd#11	1.96674e-16
C76	net31#6	y#1	8.20523e-18
C77	a#1	gnd#11	3.06374e-16
C78	y#3	vdd#14	1.92444e-17
C79	net31#2	net12#9	1.06627e-17
C80	gnd#2	net12#4	3.68329e-17
C81	b#8	vdd#50	1.97451e-16
C82	vdd#7	y#9	9.05239e-18
C83	a#1	vdd#34	1.26653e-16
C84	vdd#29	gnd#11	6.15324e-16
C85	net12#6	vdd#3	1.07589e-17
C86	gnd#13	net29	5.22889e-17
C87	y#4	net12#14	4.05599e-17
C88	net29#2	net12#10	1.93399e-18
C89	b#7	gnd#11	4.67988e-17
C90	y#8	b#6	7.39521e-18
C91	net31#3	vdd#44	3.52838e-18
C92	a#12	gnd#11	3.31852e-16
C93	net12#4	b#8	1.82453e-16
C94	net12#2	vdd#50	7.38028e-17
C95	net12	gnd#2	1.38548e-16
C96	b#1	gnd#11	3.94967e-16
C97	y#4	vdd#7	2.66547e-17
C98	y#11	vdd#22	4.19844e-17
C99	a#2	vdd#2	5.2722e-17
C100	vdd#37	a#3	1.85973e-17
C101	vdd#15	y#10	7.03723e-18
C102	net12#14	vdd#7	1.86748e-16
C103	vdd#30	gnd#11	1.00182e-16
C104	gnd#2	vdd#37	1.05786e-16
C105	gnd#10	b#7	7.09555e-18
C106	a#6	net31#3	6.36455e-17
C107	gnd#6	net12#4	8.04794e-17
C108	net12#2	gnd#11	7.0986e-17
C109	net29#2	b#6	7.73756e-19
C110	gnd#13	net29#2	1.83704e-17
C111	y#3	net12#14	7.09638e-17
C112	net12#13	net31#6	1.20562e-17
C113	vdd#37	a#12	7.37736e-17
C114	a#14	vdd#34	4.54289e-17
C115	net12#6	gnd#11	4.54162e-17
C116	vdd#50	gnd#11	3.96557e-17
C117	vdd#3	a#12	5.17623e-17
C118	vdd#31	gnd#11	1.044e-16
C119	a#6	vdd#48	3.54656e-16
C120	a#5	net31#3	4.78948e-18
C121	net12#14	vdd#5	2.81881e-17
C122	net12#11	gnd#11	9.36845e-18
C123	y#4	b#6	4.72603e-18
C124	vdd#37	a#13	9.43574e-18
C125	vdd#7	b#9	1.1592e-16
C126	vdd#50	net12#13	1.1052e-17
C127	net29#2	a#9	4.39218e-17
C128	vdd#37	a#1	1.57221e-17
C129	vdd#49	gnd#11	4.07067e-17
C130	vdd#32	gnd#11	2.23683e-16
C131	b#4	y#8	6.53797e-18
C132	vdd#7	net31	3.07312e-17
C133	net31#2	net12#12	5.91606e-18
C134	net12#15	gnd#11	2.61843e-16
C135	net12#10	net31	4.63113e-17
C136	vdd#41	gnd#11	6.24295e-17
C137	y#3	vdd#7	1.1575e-17
C138	b#8	vdd#38	2.46466e-17
C139	net31#2	gnd#11	3.37529e-17
C140	net12#6	vdd#38	6.01854e-18
C141	vdd#7	b#6	1.06075e-16
C142	net29	b#4	1.10775e-16
C143	vdd#21	gnd#11	2.40683e-16
C144	net12#9	a#5	8.34157e-18
C145	net12#4	gnd#11	1.99022e-17
C146	net31#2	vdd#47	3.96512e-17
C147	net12	b#2	1.17807e-17
C148	vdd#33	gnd#11	5.75235e-16
C149	net12#6	b#3	1.26548e-17
C150	y#3	b#6	1.33634e-17
C151	b#4	net29#2	4.89104e-17
C152	vdd#14	gnd#11	1.03101e-16
C153	y#2	vdd#7	3.45395e-17
C154	net31#6	a#5	5.0251e-18
C155	net12#14	vdd#13	5.65101e-18
C156	vdd#45	gnd#11	1.28734e-17
C157	y#8	net12#13	1.29779e-17
C158	net12#15	net28	5.26288e-17
C159	y#2	b#6	1.25274e-17
C160	net12#10	vdd#45	5.78213e-17
C161	gnd#13	b#4	1.79358e-17
C162	vdd#50	net31#6	1.77079e-17
C163	vdd#22	gnd#11	2.37921e-16
C164	a#10	y#8	5.53741e-17
C165	gnd#7	net12#15	3.7652e-17
C166	y#11	vdd#15	5.2929e-17
C167	y#8	gnd#11	9.30527e-18
C168	a#9	y#3	5.13049e-17
C169	a#5	net12#12	2.81356e-17
C170	gnd#3	a#12	6.20731e-18
C171	net12	vdd#38	9.45008e-17
C172	net12#2	vdd#37	2.59638e-17
C173	net12#4	vdd#38	1.01721e-17
C174	net28	gnd#11	9.56032e-17
C175	net28	vdd#14	8.35829e-18
C176	y#2	net31	3.1883e-16
C177	net29#2	a#10	6.92886e-17
C178	net29#2	net12#13	1.11199e-18
C179	vdd#16	b#10	2.37097e-17
C180	vdd#17	y#10	8.20864e-18
C181	net12#11	vdd#45	4.03661e-17
C182	net28#3	net12#15	1.11143e-16
C183	y#9	b#10	2.50645e-17
C184	y#12	gnd#11	1.55162e-16
C185	y#3	b#4	8.84915e-18
C186	net29	gnd#11	5.14016e-17
C187	y#3	vdd#5	3.40557e-17
C188	net12#14	gnd#11	2.05308e-16
C189	net12#10	y#1	1.53426e-16
C190	gnd#5	vdd#49	1.01094e-17
C191	b#5	net29	4.83155e-17
C192	y#3	net12#13	2.85987e-17
C193	vdd#5	net31	4.5519e-17
C194	net31#2	vdd#45	4.91607e-17
C195	y#2	vdd#5	2.19181e-16
C196	gnd#8	net28#3	1.26226e-17
C197	net29#2	gnd#11	6.87645e-17
C198	b#4	a#10	8.71314e-18
C199	net28	vdd#22	5.39096e-18
C200	net12#6	vdd#2	7.21208e-18
C201	vdd#37	gnd#11	2.06102e-16
C202	y#7	net12#14	3.76125e-17
C203	gnd#13	b#5	5.88355e-17
C204	y#12	vdd#45	3.44279e-17
C205	y#7	gnd#11	4.61701e-17
C206	net28	net12#14	5.13871e-18
C207	a#7	y#3	2.28828e-17
C208	y#2	net12#10	1.8519e-17
C209	vdd#16	gnd#11	4.27444e-17
C210	net12#13	vdd#5	1.6143e-16
C211	b#2	vdd#50	9.74644e-17
C212	a#7	b#4	1.14602e-17
C213	vdd#2	a#4	2.14827e-17
C214	b#9	gnd#11	4.5539e-17
C215	net28#3	gnd#11	5.92572e-17
C216	net12#14	vdd#14	1.57698e-17
C217	y#2	net12#9	2.84234e-17
C218	a#4	vdd#5	8.46203e-17
C219	a#7	net12#13	9.9542e-17
C220	vdd#3	gnd#11	3.40869e-17
C221	a#13	vdd#3	4.7905e-17
C222	net31#6	y#2	2.54044e-16
C223	b#10	vdd#45	2.19215e-17
C224	gnd#6	net12#3	9.11235e-17
C225	net12#10	b#6	1.65986e-17
C226	net12#4	b#2	1.69292e-16
C227	b#9	vdd#45	8.02924e-17
C228	b#6	gnd#11	1.93189e-16
C229	b#3	vdd#50	6.67376e-18
C230	vdd#5	net12#10	3.56221e-17
C231	vdd#18	gnd#11	6.57093e-17
C232	vdd#23	y#9	2.47265e-17
C233	vdd#4	y#2	7.51738e-18
C234	vdd#3	a#5	3.32337e-17
C235	net31#2	y#2	3.25633e-17
C236	a#7	vdd#5	1.45288e-16
C237	gnd#7	net28	2.05236e-17
C238	net12#10	net31#6	8.57549e-17
C239	gnd#2	vdd#38	2.90472e-17
C240	a#11	gnd#11	1.47485e-17
C241	gnd#3	a#13	3.87014e-17
C242	y#4	gnd#11	6.37126e-17
C243	a#11	vdd#41	5.13145e-17
C244	net12#14	vdd#23	6.09188e-17
C245	net12#4	vdd#50	2.23127e-16
C246	a#2	vdd#1	7.45995e-17
C247	net12	a#12	5.81571e-18
C248	b#4	net12#15	2.12432e-17
C249	a#9	gnd#11	6.31976e-17
C250	b#6	vdd#45	4.34413e-17
C251	y#2	net12#12	2.26898e-17
C252	vdd#5	net31#6	1.09358e-16
C253	vdd#4	net31	3.64489e-18
C254	net31	vdd#17	2.0615e-17
C255	vdd#4	a#6	5.44179e-17
C256	net12#14	b#9	1.91767e-17
C257	vdd#4	a#8	1.40959e-17
C258	vdd#37	gnd#1	6.61189e-17
C259	vdd#5	net12#8	7.30002e-18
C260	net31#2	vdd#48	2.07001e-17
C261	net28	y#5	1.3872e-18
C262	b#10	y#10	1.87371e-16
C263	a#9	net12#10	6.54975e-18
C264	b#7	gnd#14	5.658e-17
C265	net12#11	net31#6	2.72498e-17
C266	net12#14	b#6	5.6242e-17
C267	gnd#6	vdd#38	1.06556e-17
C268	vdd#17	b#10	2.09499e-16
C269	net12#9	vdd#45	1.77202e-17
C270	vdd#44	gnd#11	6.13269e-17
C271	y#4	vdd#23	6.4548e-17
C272	net31#3	vdd#32	4.02676e-18
C273	vdd#49	a#2	8.71855e-17
C274	b#4	gnd#11	3.71075e-16
C275	vdd#4	net31#3	1.88776e-17
C276	net12#3	gnd#14	3.34344e-17
C277	a#4	vdd#4	1.30937e-16
C278	vdd#4	a#5	1.5544e-17
C279	gnd#1	a#12	1.2008e-17
C280	net12#3	b#7	5.15296e-17
C281	gnd#5	a#13	9.13463e-18
C282	a#4	net31#6	2.47865e-17
C283	a#7	net12#8	6.09843e-17
C284	y#4	vdd#13	6.72251e-18
C285	b#4	net12#14	1.05737e-17
C286	vdd#7	gnd#11	3.51615e-17
C287	y#11	vdd#17	2.54397e-17
C288	y#12	vdd#15	8.84987e-17
C289	a#8	vdd#41	2.63735e-17
C290	gnd#10	b#3	7.49528e-18
C291	net12#3	gnd#11	7.1488e-17
C292	y#7	b#6	3.59812e-17
C293	net12#13	gnd#11	8.78323e-17
C294	y#4	net28	7.18577e-17
C295	vdd#37	gnd#5	1.70875e-17
C296	a#11	vdd#47	2.61632e-16
C297	net12#2	vdd#38	8.37827e-17
C298	vdd#22	y#12	1.60051e-16
C299	a#4	net31#2	5.73575e-17
C300	net28#3	gnd#7	5.22889e-17
C301	net31#3	vdd#47	2.97439e-16
C302	y#3	gnd#11	2.60414e-17
C303	a#7	net31#6	1.99119e-17
C304	y#3	net29	3.33219e-18
C305	net31#3	a#11	2.59556e-16
C306	a#9	b#6	8.53641e-18
C307	gnd#5	a#12	1.00916e-17
C308	vdd#34	gnd#11	4.22253e-16
C309	vdd#7	y#11	7.25332e-17
C310	a#12	vdd#49	6.81382e-18
C311	gnd#2	a#4	2.7862e-17
C312	net12#7	a#7	5.17277e-17
C313	b#9	y#10	4.0608e-17
C314	net12#12	vdd#45	1.79299e-17
C315	a#6	gnd#11	3.09869e-17
C316	net29	net12#15	5.78191e-18
C317	vdd#37	b#8	5.93711e-18
C318	a#4	vdd#50	7.45917e-18
C319	vdd#40	gnd#11	1.90921e-17
C320	vdd#23	b#9	2.16977e-17
C321	vdd#23	gnd#11	5.93121e-17
C322	vdd#3	net31#6	8.39304e-18
C323	vdd#2	a#6	1.60407e-17
C324	vdd#50	net29#2	7.35582e-18
C325	a#6	vdd#41	6.19438e-17
C326	a#1	vdd#49	1.3311e-17
C327	net28#3	y#5	2.47647e-18
C328	net12#9	net31	2.14091e-16
C329	net31#2	vdd#44	2.6693e-17
C330	gnd#2	a#7	3.4007e-17
C331	net12#3	b#2	1.92673e-17
C332	y#9	vdd#21	1.97221e-17
C333	vdd#4	net31#6	7.38357e-18
C334	b#9	vdd#17	3.5607e-16
C335	a#5	gnd#11	2.32252e-16
C336	gnd#14	b#3	2.80066e-17
C337	net12#2	b#8	1.12609e-17
C338	y#1	net12#9	1.87374e-16
C339	a#9	net12#13	6.73114e-17
C340	a#7	vdd#50	4.85567e-17
C341	net28#3	y#4	1.86963e-17
C342	vdd#5	gnd#11	4.20109e-17
C343	vdd#22	y#9	5.84091e-18
C344	gnd#6	a#7	8.93465e-18
C345	gnd#6	b#2	2.46438e-17
C346	vdd#14	avC10	4.06992e-18
C347	vdd#6	net31#3	3.55036e-18
C348	y#10	avC10	4.75715e-16
C349	vdd#6	net31	1.06579e-17
C350	avC10	vdd#45	5.58308e-17
C351	vdd#7	avC10	2.98549e-18
C352	b#10	avC10	2.17277e-17
C353	vdd#16	avC10	2.13559e-17
C354	vdd#17	avC10	2.4857e-18
C355	vdd#6	net31#2	1.5482e-17
C356	vdd#23	avC10	5.64619e-17
C357	avC10	vdd#20	4.97058e-18
C358	vdd#15	avC10	5.59875e-16
C359	y#9	avC10	6.96952e-16
C360	vdd#22	avC10	2.71428e-17
C361	vdd#6	y#9	2.78454e-17
C362	b#9	avC10	2.41482e-17
C363	a#11	vdd#6	1.40223e-17
C364	vdd#6	gnd#11	1.40159e-16
C365	vdd#38	gnd#11	5.83761e-18
C366	gnd#2	vdd#3	7.73588e-18
C367	vdd#4	a#2	1.24695e-18
C368	vdd#1	a#6	1.41785e-18
C369	vdd#2	a#5	1.45616e-18
C370	vdd#44	a#5	1.78429e-18
C371	a#12	vdd#1	2.93045e-18
C372	vdd#50	a#12	3.14103e-18
C373	vdd#50	a#13	3.21557e-18
C374	vdd#48	a#5	3.26347e-18
C375	a#4	vdd#45	3.32852e-18
C376	vdd#2	a#14	3.51987e-18
C377	vdd#50	a#3	3.65044e-18
C378	vdd	a#11	4.06662e-18
C379	vdd#2	a#12	4.14661e-18
C380	vdd#47	a#8	4.21227e-18
C381	vdd#44	a#11	4.67732e-18
C382	vdd#32	a#8	4.69152e-18
C383	vdd#33	a#14	4.69152e-18
C384	vdd#5	a#9	4.818e-18
C385	vdd#48	a#11	5.46805e-18
C386	b#10	vdd#26	2.00114e-18
C387	vdd#14	b#6	2.77783e-18
C388	vdd#23	b#6	3.23648e-18
C389	vdd#14	b#9	3.5182e-18
C390	vdd#5	b#6	4.30759e-18
C391	a#4	gnd#5	2.73698e-18
C392	gnd#2	a#12	5.67837e-18
C393	y#11	vdd#18	1.00637e-18
C394	vdd#16	y#10	1.02354e-18
C395	y#10	vdd#20	1.07484e-18
C396	vdd#5	y#1	1.26184e-18
C397	y#11	vdd#21	1.75003e-18
C398	vdd#23	y#5	1.78368e-18
C399	vdd#6	y#2	1.91786e-18
C400	vdd#6	y#11	2.3985e-18
C401	vdd#23	y#10	2.45644e-18
C402	vdd#14	y#5	2.7492e-18
C403	vdd#7	y#7	2.81704e-18
C404	vdd#14	y#10	3.14e-18
C405	y#4	vdd#45	3.21568e-18
C406	y#2	vdd#17	3.93003e-18
C407	y#2	vdd#45	4.70219e-18
C408	y#12	vdd#21	5.10537e-18
C409	y#12	vdd#18	5.49479e-18
C410	gnd#14	b#2	1.62737e-18
C411	gnd#9	b#5	1.77961e-18
C412	a#7	b#6	1.76924e-18
C413	a#10	b#6	3.02715e-18
C414	vdd#3	net31#2	2.08592e-18
C415	net31#3	vdd#41	2.38984e-18
C416	vdd#7	net31#6	2.66951e-18
C417	net31#2	vdd#41	3.19696e-18
C418	vdd#17	net12#9	1.39539e-18
C419	vdd#50	net12#11	1.79785e-18
C420	net12#15	vdd#14	2.609e-18
C421	net12#6	vdd#7	3.7037e-18
C422	vdd#50	net12#8	3.74732e-18
C423	net12	vdd#49	3.87378e-18
C424	net12	vdd#37	4.40638e-18
C425	vdd#5	net12#11	5.00291e-18
C426	net12#15	vdd#13	5.50593e-18
C427	y#1	a#5	3.57546e-18
C428	y#2	a#9	3.6099e-18
C429	y#2	a#5	4.24114e-18
C430	y#7	b#4	3.93959e-18
C431	y#11	b#9	4.17098e-18
C432	y#9	b#9	4.39429e-18
C433	gnd#2	net12#6	2.96134e-18
C434	gnd#8	net12#15	3.39295e-18
C435	gnd#2	net12#13	3.88796e-18
C436	gnd#8	net12#16	4.15259e-18
C437	net12#6	gnd#14	4.91746e-18
C438	gnd#10	net12#3	5.05022e-18
C439	y#4	avC10	1.55645e-18
C440	net12#6	a#5	2.00943e-18
C441	a#7	net12#11	2.26815e-18
C442	a#7	net12#4	4.24794e-18
C443	net31	b#9	1.64513e-18
C444	b#8	net12#13	1.03511e-18
C445	net12#4	b#3	1.12264e-18
C446	net12#8	b#6	1.57256e-18
C447	net12	b#8	1.66749e-18
C448	net12#2	b#2	1.76957e-18
C449	net12#6	b#2	1.9458e-18
C450	net12#6	b#8	2.57585e-18
C451	net31#2	y#1	2.92761e-18
C452	y#8	net12#10	2.4355e-18
C453	y#2	net12#13	2.61815e-18
C454	net12#15	y#5	2.67103e-18
C455	y#2	net12#8	3.07359e-18
C456	net12#14	y#5	5.28842e-18
C457	net12#6	y#2	5.54093e-18
C458	net31#6	net12#9	2.56038e-18
C459	net31	net12#12	2.5699e-18
C460	avC10	gnd	6.81928e-18
C461	b#10	gnd	4.37385e-18
C462	a#11	gnd	1.80265e-18
C463	net12#9	gnd	8.94911e-19
C464	net12#12	gnd	1.05737e-18
C465	b#8	gnd	5.22198e-18
C466	vdd#13	gnd	4.63783e-21
C467	a#10	gnd	1.31675e-20
C468	b#5	gnd	2.32469e-18
C469	a#13	gnd	2.13953e-18
C470	b#7	gnd	1.60778e-18
C471	vdd#20	gnd	8.54884e-19
C472	net12#15	gnd	1.00252e-19
C473	vdd#14	gnd	1.33559e-18
C474	vdd#8	gnd	5.18559e-19
C475	net12#14	gnd	1.92882e-18
C476	b#9	gnd	4.10276e-18
C477	b#6	gnd	2.46163e-18
C478	a#9	gnd	5.0824e-18
C479	b#4	gnd	1.08236e-17
C480	net12#13	gnd	6.03614e-19
C481	a#6	gnd	1.23151e-18
C482	a#5	gnd	1.24152e-17
C483	net12#8	gnd	9.6565e-19
C484	b#3	gnd	3.91708e-19
C485	a#2	gnd	2.83814e-18
C486	a#3	gnd	3.43291e-18
C487	a#1	gnd	5.43706e-19
C488	net12#6	gnd	8.23524e-18
C489	net12	gnd	6.21231e-18
C490	vdd#21	gnd	1.01483e-18
C491	y#12	gnd	8.43516e-19
C492	vdd#12	gnd	1.01506e-19
C493	vdd#16	gnd	1.33133e-18
C494	y#9	gnd	2.97443e-18
C495	y#4	gnd	2.45666e-18
C496	vdd#6	gnd	3.18386e-18
C497	vdd#7	gnd	3.87477e-19
C498	y#3	gnd	1.48759e-18
C499	y#2	gnd	2.19189e-18
C500	vdd#5	gnd	5.75101e-19
C501	a#4	gnd	1.54121e-18
C502	a#7	gnd	3.04878e-18
C503	vdd#4	gnd	7.28726e-19
C504	net12#7	gnd	1.18772e-18
C505	net12#2	gnd	8.06591e-19
C506	vdd#41	gnd	1.23185e-18
C507	vdd#45	gnd	1.2367e-18
C508	net28	gnd	4.36406e-18
C509	y#5	gnd	5.19824e-19
C510	net28#3	gnd	5.66865e-18
C511	vdd#15	gnd	2.60124e-18
C512	y#10	gnd	5.18559e-19
C513	vdd#40	gnd	1.19699e-18
C514	vdd#17	gnd	1.65577e-18
C515	vdd#47	gnd	8.32169e-19
C516	net31	gnd	4.83864e-18
C517	net31#3	gnd	1.70338e-18
C518	net31#6	gnd	3.91845e-18
C519	vdd#1	gnd	6.29932e-19
C520	vdd#50	gnd	2.79389e-19
C521	vdd#49	gnd	2.97698e-18
C522	net12#4	gnd	1.22635e-18
C523	y#8	gnd	1.3648e-18
C524	net29	gnd	1.26226e-17
C525	net29#2	gnd	1.00252e-19
C526	vdd#3	gnd	1.1406e-18
C527	vdd#34	gnd	3.08516e-19
C528	vdd#2	gnd	3.02635e-19
C529	net12#10	gnd	2.40707e-18
C530	net12#11	gnd	1.13345e-18
C531	net31#2	gnd	6.09218e-19
C532	y#7	gnd	4.76388e-18
C533	y#11	gnd	6.18767e-18
C534	vdd#23	gnd	6.32766e-19
C535	vdd#26	gnd	6.0577e-20
C536	vdd#31	gnd	6.05667e-19
C537	vdd#37	gnd	5.37031e-18
C538	vdd#44	gnd	9.65952e-19
*
*
.ENDS XOR2X1
*
