*
*
*
*                       LINUX           Tue May 25 13:33:05 2021
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus - (64-bit)
*  Version        : 20.1.1-s233
*  Build Date     : Wed Mar 25 13:13:47 PDT 2020
*
*  HSPICE LIBRARY
*
*
*
.GLOBAL vdd gnd
*
.SUBCKT XOR2X1 a b y
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
M6	net29#2	b#12	gnd	gnd	N_18_MM	L=1.8e-07
+ W=4.8e-07	effW=4.8e-07
M7	net28	net12#12	gnd	gnd	N_18_MM	L=1.8e-07
+ W=4.8e-07	effW=4.8e-07
M9	net11#3	a#9	gnd	gnd	N_18_MM	L=1.8e-07
+ W=2.4e-07	effW=2.4e-07
M10	net12#5	b#9	gnd	gnd	N_18_MM	L=1.8e-07
+ W=2.4e-07	effW=2.4e-07
M4	y#7	a#6	net29	gnd	N_18_MM	L=1.8e-07
+ W=4.8e-07	effW=4.8e-07
M5	y#3	net11#11	net28#4	gnd	N_18_MM
+ L=1.8e-07	W=4.8e-07
+ effW=4.8e-07
M3	y#1	b#16	net30#4	vdd	P_18_MM	L=1.8e-07
+ W=6.36e-06	effW=6.36e-06
M2	y#8	net12#10	net31#4	vdd	P_18_MM
+ L=1.8e-07	W=6.36e-06
+ effW=6.36e-06
M11	net12#2	b#8	vdd	vdd	P_18_MM	L=1.8e-07
+ W=3.18e-06	effW=3.18e-06
M0	net31	a#8	vdd	vdd	P_18_MM	L=1.8e-07
+ W=6.36e-06	effW=6.36e-06
M8	net11	a#10	vdd	vdd	P_18_MM	L=1.8e-07
+ W=3.18e-06	effW=3.18e-06
M1	net30	net11#9	vdd	vdd	P_18_MM	L=1.8e-07
+ W=6.36e-06	effW=6.36e-06
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rh1	b#8	b#4	   85.1145	$PLY_C
Rh2	b#9	b#6	   27.8221	$PLY_C
Rh3	b#6	b#10	   30.4206	$PLY_C
Rh4	b#10	b#11	   86.3343	$PLY_C
Rh5	b#11	b#2	   21.2243	$PLY_C
Rh6	b#10	b#3	  110.3262	$PLY_C
Rh7	b#11	b#5	   39.0050	$PLY_C
Rh8	b#5	b#12	   23.8666	$PLY_C
Rh9	net12#10	net12#9	  154.4446	$PLY_C
Rh10	net12#9	net12#11	   93.4606	$PLY_C
Rh11	net12#11	net12	   55.4494	$PLY_C
Rh12	net12	net12#12	   23.6444	$PLY_C
Rh13	net12#11	net12#4	  103.6595	$PLY_C
Rh14	a#6	a#5	   24.2347	$PLY_C
Rh15	a#5	a#4	  436.4613	$PLY_C
Rh16	a#4	a#7	   81.3616	$PLY_C
Rh17	a#7	a#3	  164.7824	$PLY_C
Rh18	a#3	a#1	   38.4487	$PLY_C
Rh19	a#4	a#8	  154.4884	$PLY_C
Rh20	a#7	a#9	  160.0426	$PLY_C
Rh22	a#3	a#10	   84.2131	$PLY_C
Rh23	net11#9	net11#7	  158.1077	$PLY_C
Rh24	net11#7	net11#10	  143.7236	$PLY_C
Rh25	net11#10	net11#5	   35.8910	$PLY_C
Rh26	net11#10	net11#8	  287.5862	$PLY_C
Rh27	net11#8	net11#11	   27.0923	$PLY_C
Rh28	b#16	b#13	  154.6152	$PLY_C
Rh29	b#13	b#14	   32.9050	$PLY_C
Rg1	b	b#1	    1.5566	$ME1_C
Rg2	b#1	b#2	   12.0000	$ME1_C
Rg3	a	a#1	   13.9558	$ME1_C
Rg4	b#3	b#4	   24.2543	$ME1_C
Rg5	net11	net11#2	    9.2209	$ME1_C
Rg6	net12#2	net12#3	    9.2201	$ME1_C
Rg7	net12#4	net12#6	   12.2306	$ME1_C
Rg8	net12#6	net12#7	3.881e-03	$ME1_C
Rg9	net12#6	net12#8	3.082e-02	$ME1_C
Rg10	net12#5	net12#6	   15.0000	$ME1_C
Rg11	net12#5	net12#7	   15.0000	$ME1_C
Rg12	net11#3	net11#4	   21.9633	$ME1_C
Rg13	net29	net29#2	   31.2855	$ME1_C
Rg14	net31	net31#2	    1.8788	$ME1_C
Rg15	net31#2	net31#3	1.941e-03	$ME1_C
Rg16	net31#3	net31#4	    2.4835	$ME1_C
Rg17	net31	net31#2	   15.0000	$ME1_C
Rg18	net31	net31#3	   15.0000	$ME1_C
Rg19	net28	net28#2	   15.0214	$ME1_C
Rg20	net28#2	net28#3	    7.7046	$ME1_C
Rg21	net28	net28#2	   15.0000	$ME1_C
Rg22	net11#5	net11#6	   18.5000	$ME1_C
Rg23	net28#4	net28#5	   21.6739	$ME1_C
Rg24	net30	net30#2	    1.8788	$ME1_C
Rg25	net30#2	net30#3	1.941e-03	$ME1_C
Rg26	net30#3	net30#4	    2.4841	$ME1_C
Rg27	net30	net30#2	   15.0000	$ME1_C
Rg28	net30	net30#3	   15.0000	$ME1_C
Rg29	b#14	b#15	   18.6257	$ME1_C
Rg30	y	y#2	    2.8068	$ME1_C
Rg31	y#2	y#4	    2.0124	$ME1_C
Rg32	y#4	y#5	1.691e-02	$ME1_C
Rg33	y#5	y#6	    0.9682	$ME1_C
Rg34	y#6	y#7	   15.1486	$ME1_C
Rg35	y#6	y#8	    2.5339	$ME1_C
Rg36	y#1	y#2	    1.1538	$ME1_C
Rg37	y#3	y#4	   15.0000	$ME1_C
Rg38	y#3	y#5	   15.0000	$ME1_C
Rf1	b#1	b#7	   13.0000	$ME2_C
Rf2	net12#3	net12#8	    7.3347	$ME2_C
Rf3	net11#6	net11#4	    0.5242	$ME2_C
Rf4	net11#4	net11#2	    1.7578	$ME2_C
Rf5	net28#5	net28#3	    0.3937	$ME2_C
Rf6	b#17	b#15	    6.8699	$ME2_C
Re1	b#17	b#7	    1.9800	$ME3_C
*
*       CAPACITOR CARDS
*
*
C1	net28#5	a#6	2.9326e-18
C2	net12#10	y#8	4.1633e-16
C3	b#17	y#3	9.2882e-18
C4	net12#9	y#8	1.22467e-16
C5	net12#8	b#6	1.80862e-17
C6	net11#9	vdd	4.61606e-16
C7	b#16	vdd	1.42804e-17
C8	net12#3	b#8	2.47541e-17
C9	a#8	vdd	4.76103e-16
C10	a#4	net11#5	3.1261e-17
C11	net12#10	vdd	1.5361e-17
C12	a#10	vdd	2.30786e-16
C13	net11#6	net31	4.75902e-18
C14	net31#4	net12#10	3.73894e-16
C15	a#5	net12#9	1.03555e-16
C16	b#8	vdd	2.18135e-16
C17	b#14	vdd	3.02613e-17
C18	net11#10	net30#4	4.90006e-16
C19	b#13	vdd	2.58192e-17
C20	net12#5	net11#3	8.24944e-18
C21	net11#8	vdd	9.75624e-17
C22	net11#7	vdd	3.14695e-16
C23	a#5	vdd	2.01207e-16
C24	net12#9	vdd	4.23635e-17
C25	net31	a#4	2.82717e-16
C26	a#4	vdd	4.82256e-16
C27	a#3	vdd	3.89356e-16
C28	net12#9	net31#4	1.47084e-16
C29	b#4	vdd	1.35224e-16
C30	b#3	vdd	6.43933e-17
C31	net28#3	a#6	1.33497e-17
C32	a#1	vdd	2.15682e-16
C33	b#17	vdd	3.80646e-17
C34	b#7	vdd	1.48086e-17
C35	b#17	net28#4	2.28598e-18
C36	net11#6	vdd	9.4479e-18
C37	net31	a#7	3.79651e-18
C38	net11#4	vdd	1.42397e-16
C39	net28	net12#11	7.63393e-18
C40	net11#2	vdd	7.06312e-16
C41	net12#3	vdd	4.32915e-16
C42	net30	vdd	1.01929e-15
C43	y#1	vdd	1.86059e-16
C44	net31	vdd	7.57646e-16
C45	vdd	net31#4	5.50035e-18
C46	net11	vdd	2.69836e-17
C47	vdd	net12#2	1.37036e-17
C48	y#8	a#4	3.2348e-16
C49	net11#6	y#8	7.77297e-17
C50	net29#2	vdd	1.57154e-17
C51	a#7	vdd	2.50359e-16
C52	net11#10	vdd	2.61755e-16
C53	y#6	vdd	8.31636e-18
C54	net28	net29	1.40673e-17
C55	y#6	net28#4	6.27456e-18
C56	a#10	net11	1.61578e-16
C57	net31#4	a#4	5.91991e-18
C58	b#17	y#6	1.77951e-17
C59	y#7	a#5	1.71041e-17
C60	b#15	y#3	1.28598e-16
C61	net11#4	net31	4.75442e-17
C62	net12#11	net31#4	3.74218e-18
C63	net12#4	net31#4	2.33448e-17
C64	net29	a#5	6.15161e-17
C65	net29#2	net12#5	1.2979e-18
C66	net11#10	b#16	6.13955e-17
C67	b#8	net12#2	1.61579e-16
C68	net11#4	y#8	2.03714e-17
C69	y#8	net11#10	1.55952e-17
C70	b#17	net28#5	1.79441e-17
C71	y#3	net28#5	1.21628e-17
C72	b#7	net29	3.35923e-18
C73	net29	net12#9	7.07609e-17
C74	net11#4	net31#4	1.27234e-16
C75	b#17	net11#6	2.91866e-17
C76	net12#3	b#4	3.23379e-17
C77	net12#8	y#8	6.67626e-18
C78	b#17	net11#8	1.34576e-17
C79	net11#2	net31	2.31503e-17
C80	a#3	net11	1.00075e-16
C81	net11#11	y#3	6.92895e-17
C82	net29	y#6	1.10153e-17
C83	net28#4	net11#11	4.82104e-17
C84	b#17	net28#3	1.57332e-17
C85	net12#2	a#3	4.71822e-18
C86	net28#5	y#7	1.48703e-18
C87	net12#3	b#3	4.38566e-18
C88	net12#8	net31#4	2.33762e-17
C89	net28	net29#2	8.99893e-18
C90	net11#2	a#1	8.43471e-18
C91	net12#3	net31	5.28287e-18
C92	b#5	net12#4	3.64001e-17
C93	net29	net31#4	1.83004e-17
C94	y#1	net30	1.11399e-16
C95	net29#2	net12#9	1.41807e-17
C96	net28#5	net11#8	1.07764e-17
C97	net28#5	net29	2.60322e-18
C98	b#7	net29#2	3.62555e-17
C99	b#6	net31#4	6.83705e-18
C100	a#6	y#7	4.79082e-17
C101	net11#7	b#16	1.75505e-17
C102	y#6	net30#4	1.38611e-17
C103	net12#2	a#7	1.71537e-16
C104	b#7	net11#4	3.12998e-17
C105	net29	a#6	4.83619e-17
C106	b#7	net28	9.93904e-18
C107	b#17	a#5	7.3223e-18
C108	b#4	a#7	2.94966e-17
C109	net28#5	y#6	1.06645e-16
C110	y#3	net28#4	1.04912e-16
C111	b#5	net31#4	9.42148e-18
C112	y#6	b#13	1.28794e-17
C113	net12#3	net31#4	6.62302e-18
C114	b#7	net12#8	1.31428e-17
C115	net28#3	y#7	6.44039e-17
C116	net30#4	y#1	5.36459e-16
C117	net12#5	net31#4	1.39209e-17
C118	net12#10	a#5	2.06125e-17
C119	b#7	net12#9	4.70554e-18
C120	net29#2	net12#4	2.14448e-17
C121	b#14	y#1	7.14738e-17
C122	net28#3	net29	9.96084e-17
C123	b#8	a#7	2.64412e-17
C124	y#8	net30	9.20487e-18
C125	net12#10	a#4	6.1857e-17
C126	net29#2	net31#4	7.13656e-17
C127	y#6	net11#8	2.9407e-17
C128	net12	b#5	5.30416e-18
C129	b#7	net12#3	7.05096e-18
C130	b#13	y#1	1.3797e-16
C131	net28#3	a#5	1.04134e-17
C132	net29#2	y#6	3.86281e-18
C133	net12#3	a#7	3.31412e-17
C134	b#17	net30	3.88665e-18
C135	b#13	net30#4	1.37547e-16
C136	b#7	net12#4	1.40803e-17
C137	b#9	net12#5	4.53375e-17
C138	b#11	net12#4	7.39526e-18
C139	net28#3	y#6	6.6572e-17
C140	a#5	net11#10	1.4911e-17
C141	b#8	a#3	2.35784e-17
C142	b#17	y#1	8.12749e-17
C143	net11#6	a#4	8.59904e-18
C144	b#4	net12#2	7.52761e-17
C145	y#8	net30#4	7.39757e-17
C146	net11#8	net30#4	1.62332e-16
C147	net11#7	net30	2.57337e-16
C148	net29	net12#11	5.28951e-18
C149	b#17	net30#4	3.51695e-17
C150	net12#5	b#6	8.48578e-18
C151	net31#4	y#6	4.06672e-17
C152	y#3	b#14	2.93036e-17
C153	net29	y#7	4.12117e-17
C154	b#12	net29#2	5.376e-17
C155	net12#8	net11#3	1.57804e-17
C156	net31	y#8	1.12041e-16
C157	net11#4	a#4	4.05688e-17
C158	net11#9	net30	3.86783e-16
C159	net12#8	net11#4	8.67288e-18
C160	net11#8	b#13	1.05666e-16
C161	net31	net11#7	6.13756e-18
C162	net12	net29	1.85766e-17
C163	b#15	y#1	6.35592e-17
C164	y#3	b#13	1.11292e-17
C165	b#9	net12#4	9.6612e-18
C166	b#17	y#8	2.64111e-17
C167	net30	b#16	1.87245e-17
C168	net28#4	b#13	1.66351e-18
C169	b#16	y#1	4.14391e-16
C170	net29#2	b#5	2.9207e-17
C171	net12#12	net28	5.06872e-17
C172	a#4	net11#10	2.36792e-17
C173	net30#4	b#16	3.77531e-16
C174	net30	net11#10	9.32351e-18
C175	net12#8	net29#2	3.24014e-18
C176	y#6	a#5	1.01066e-16
C177	y#3	net11#8	3.99278e-17
C178	net30#4	a#5	1.09593e-17
C179	net12#3	net11#4	9.08697e-17
C180	net31#4	y#8	4.85173e-16
C181	a#5	net11#8	2.00549e-17
C182	net12#3	net11#3	2.26579e-17
C183	net28#4	net11#8	1.93836e-17
C184	net12	net29#2	1.4044e-17
C185	a#8	net31	3.9043e-16
C186	b#7	net31#4	2.86246e-17
C187	net30	a#4	4.12897e-18
C188	a#3	net11#2	3.58884e-17
C189	net11#2	a#10	2.69289e-17
C190	a#5	y#8	3.42398e-16
C191	net28#5	net11#11	2.90522e-18
C192	net28	net12	4.93419e-17
C193	b#1	net12#4	4.20742e-18
C194	net12#9	y#6	3.48683e-17
C195	net12	b#12	8.8627e-18
C196	b#12	net12#11	1.33088e-17
C197	net12#8	b#10	5.84843e-18
C198	net11#6	net30#4	2.74706e-17
C199	net29#2	net12#11	1.25345e-16
C200	net12#3	a#3	1.53228e-17
C201	a#4	net11#7	1.43409e-17
C202	net31	net12#10	1.52962e-17
C203	net12#3	net11#2	2.41171e-17
C204	net28#4	net30#4	1.1344e-17
C205	net30#4	a#4	7.28985e-18
C206	a#9	b#4	3.10026e-17
C207	a#9	net12#3	1.10519e-17
C208	b#10	a#9	1.93338e-17
C209	b#6	a#9	5.23298e-17
C210	net11#4	a#9	6.46015e-18
C211	a#9	net31#4	1.30013e-17
C212	b#3	a#9	1.67447e-17
C213	net11#3	a#9	1.76545e-16
C214	net12#8	a#9	1.74404e-17
C215	net11#3	net12#2	1.56395e-18
C216	net11#3	net12#4	2.8902e-18
C217	net11#4	net12#10	4.0643e-18
C218	net30#4	net11#7	3.729e-18
C219	a#9	net12#10	1.44633e-18
C220	net12	a#5	1.76204e-18
C221	a#9	net12#2	3.75151e-18
C222	net31#4	a#5	2.52419e-18
C223	b#17	net11#10	2.05208e-18
C224	b#17	net11#4	2.34034e-18
C225	b#15	net11#8	2.50862e-18
C226	b#7	net11#3	3.95347e-18
C227	net11#4	b#4	5.15305e-18
C228	b#7	net12#11	1.97449e-18
C229	b#17	net12#9	2.23396e-18
C230	b#7	net12#10	2.29194e-18
C231	b#7	net12	2.65937e-18
C232	b#5	net12#11	3.13329e-18
C233	net11#6	y#1	3.29572e-18
C234	y#8	net11#8	3.59261e-18
C235	y#8	net11#5	4.18539e-18
C236	y#1	net11#10	4.30986e-18
C237	b#4	net31	2.15858e-18
C238	b#17	net31	2.92132e-18
C239	net28#3	net12#9	1.10418e-18
C240	vdd	gnd	2.24966e-15
C241	a	gnd	3.12656e-16
C242	b	gnd	2.39349e-16
C243	y	gnd	4.37546e-16
C244	b#16	gnd	7.14811e-19
C245	a#8	gnd	1.16897e-18
C246	net12#10	gnd	2.46514e-18
C247	b#8	gnd	1.33416e-18
C248	net11#11	gnd	3.04321e-17
C249	a#6	gnd	5.21299e-17
C250	a#9	gnd	3.34079e-16
C251	b#9	gnd	8.54491e-17
C252	b#12	gnd	7.27594e-17
C253	net12#12	gnd	9.64534e-17
C254	b#14	gnd	6.32309e-17
C255	b#13	gnd	3.3736e-17
C256	net11#8	gnd	1.42668e-16
C257	net11#7	gnd	9.6234e-17
C258	net11#5	gnd	1.18391e-16
C259	a#5	gnd	1.2481e-16
C260	net12#9	gnd	5.04387e-17
C261	a#4	gnd	1.25317e-16
C262	net12#4	gnd	1.32071e-16
C263	a#3	gnd	9.16258e-17
C264	b#6	gnd	1.96369e-16
C265	b#5	gnd	2.40818e-16
C266	net12	gnd	2.95787e-16
C267	b#4	gnd	3.53062e-17
C268	b#3	gnd	2.20083e-16
C269	a#1	gnd	3.24547e-16
C270	b#2	gnd	9.71299e-17
C271	b#17	gnd	1.4218e-16
C272	b#7	gnd	1.78722e-16
C273	b#15	gnd	3.67068e-17
C274	net28#5	gnd	9.03856e-17
C275	net11#6	gnd	8.50665e-17
C276	net28#3	gnd	2.16589e-16
C277	net11#4	gnd	8.04669e-17
C278	net12#8	gnd	6.65289e-17
C279	net11#2	gnd	4.53506e-17
C280	net12#3	gnd	2.28237e-17
C281	b#1	gnd	2.91157e-16
C282	net30	gnd	3.79168e-17
C283	y#1	gnd	3.01254e-16
C284	net30#4	gnd	6.28199e-18
C285	net31	gnd	2.3352e-17
C286	y#8	gnd	2.08094e-18
C287	net31#4	gnd	6.7061e-18
C288	net11	gnd	1.40348e-18
C289	net12#2	gnd	1.06289e-18
C290	y#3	gnd	3.95166e-16
C291	net28#4	gnd	5.39924e-18
C292	y#7	gnd	4.53272e-18
C293	net29	gnd	7.42985e-17
C294	net11#3	gnd	6.34246e-17
C295	net12#5	gnd	7.65625e-17
C296	net29#2	gnd	1.13421e-16
C297	net28	gnd	2.55625e-16
C298	b#10	gnd	2.76132e-16
C299	b#11	gnd	1.57694e-16
C300	net12#11	gnd	2.03726e-16
C301	a#7	gnd	7.6762e-17
C302	net11#10	gnd	2.08472e-17
C303	y#6	gnd	1.46049e-16
*
*
.ENDS XOR2X1
*
