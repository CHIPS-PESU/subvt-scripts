*
*
*
*                       LINUX           Tue May 18 23:29:22 2021
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus - (64-bit)
*  Version        : 20.1.1-s233
*  Build Date     : Wed Mar 25 13:13:47 PDT 2020
*
*  HSPICE LIBRARY
*
*
*

*
.SUBCKT XNOR2X1 gnd b y
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
M9	avC3#13	avC3#47	gnd#3	gnd#13	n_18_mm
+ L=1.8e-07	W=2.4e-07
+ effW=2.4e-07
M10	net037	b#10	gnd#9	gnd#13	n_18_mm	L=1.8e-07
+ W=2.4e-07	effW=2.4e-07
M4	y#8	avC3#46	net017#2	gnd#13	n_18_mm
+ L=1.8e-07	W=4.8e-07
+ effW=4.8e-07
M6	net017	net037#12	gnd#11	gnd#13	n_18_mm
+ L=1.8e-07	W=4.8e-07
+ effW=4.8e-07
M5	y#10	avC3#37	net013#5	gnd#13	n_18_mm
+ L=1.8e-07	W=4.8e-07
+ effW=4.8e-07
M7	net013	b#14	gnd#7	gnd#13	n_18_mm	L=1.8e-07
+ W=4.8e-07	effW=4.8e-07
M8	avC3#11	avC3#48	avC10	avC3#65	p_18_mm
+ L=1.8e-07	W=3.18e-06
+ effW=3.18e-06
M11	net037#5	b#11	avC5	avC3	p_18_mm	L=1.8e-07
+ W=3.18e-06	effW=3.18e-06
MavD28_3_unmatched	y#1	avS52	avC3#64	avC3#61	p_18_mm
+ L=1.8e-07	W=3.18e-06
+ effW=3.18e-06
MavD28_4_unmatched	avC3#57	avC3#17	avC3#63	avC3#53
+ p_18_mm	L=1.8982e-07	W=3.31e-06	effW=3.31e-06
MavD28_5_unmatched	avC9	avC3#52	avC3#57	avC3#53
+ p_18_mm	L=1.8e-07	W=3.18e-06	effW=3.18e-06
MavD28_6_unmatched	avC3#21	b#5	y#1	avC3#61	p_18_mm
+ L=1.8e-07	W=3.18e-06
+ effW=3.18e-06
MavD28_7_unmatched	y#4	avS50	avC3#41	avC3#61	p_18_mm
+ L=1.8e-07	W=3.18e-06
+ effW=3.18e-06
MavD28_8_unmatched	avC3#33	avC3#51	avC8	avC3#53
+ p_18_mm	L=1.8207e-07	W=3.3175e-06	effW=3.3175e-06
MavD28_9_unmatched	avC3#40	net037#10	y#4	avC3#61
+ p_18_mm	L=1.8e-07	W=3.18e-06	effW=3.18e-06
MavD28_10_unmatched	avC7	avC3#43	avC3#33	avC3#53
+ p_18_mm	L=1.8196e-07	W=3.31e-06	effW=3.31e-06
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rh1	avC3#17	avC3#16	   78.4924	$PLY_C
Rh2	b#5	b#6	  170.1728	$PLY_C
Rh3	b#6	b#7	   95.8988	$PLY_C
Rh4	b#7	b#3	   93.5989	$PLY_C
Rh5	b#3	b#2	   25.0791	$PLY_C
Rh6	b#2	b#8	    2.6059	$PLY_C
Rh7	b#8	b#1	   65.5443	$PLY_C
Rh9	b#7	b#9	  130.9705	$PLY_C
Rh10	b#3	b#10	   28.7860	$PLY_C
Rh11	b#8	b#11	   82.8780	$PLY_C
Rh12	avC3#37	avC3#31	   23.4666	$PLY_C
Rh13	avC3#31	avC3#23	   32.4036	$PLY_C
Rh14	b#14	b#13	   23.4666	$PLY_C
Rh15	b#13	b#12	   32.4036	$PLY_C
Rh16	net037#10	net037#11	  173.0526	$PLY_C
Rh17	net037#11	net037#8	  265.7966	$PLY_C
Rh19	net037#8	net037#12	   23.6035	$PLY_C
Rh20	net037#8	net037#4	  233.3419	$PLY_C
Rh21	avC3#43	avC3#39	   69.4665	$PLY_C
Rh22	avC3#39	avC3#44	  212.2646	$PLY_C
Rh23	avC3#44	avC3#10	  133.1560	$PLY_C
Rh24	avC3#10	avC3#7	   93.0094	$PLY_C
Rh26	avC3#39	avC3#45	   16.2206	$PLY_C
Rh27	avC3#45	avC3#42	   33.7109	$PLY_C
Rh28	avC3#44	avC3#19	  298.6376	$PLY_C
Rh29	avC3#19	avC3#46	   24.4031	$PLY_C
Rh30	avC3#7	avC3#8	   23.5153	$PLY_C
Rh31	avC3#8	avC3#47	   27.4073	$PLY_C
Rh32	avC3#7	avC3#48	   84.1337	$PLY_C
Rh33	avC3#45	avC3#49	    0.3081	$PLY_C
Rh34	avC3#49	avC3#50	    1.0406	$PLY_C
Rh35	avC3#50	avC3#51	   66.3792	$PLY_C
Rh36	avC3#42	avC3#52	  141.7952	$PLY_C
Rh37	avC3#27	avC3#45	   12.0000	$PLY_C
Rh38	avC3#30	avC3#49	   12.0000	$PLY_C
Rh39	avC3#32	avC3#50	   12.0000	$PLY_C
Rg2	avC3#2	avC3#4	    6.6851	$ME1_C
Rg3	avC3	avC3#2	   15.0000	$ME1_C
Rg4	avC3	avC3#2	   15.0000	$ME1_C
Rg5	b#1	b	   13.3849	$ME1_C
Rg6	gnd#1	gnd#3	   16.2850	$ME1_C
Rg7	net037#2	net037#3	5.094e-03	$ME1_C
Rg8	net037#3	net037#4	   12.1809	$ME1_C
Rg9	net037	net037#2	   15.0000	$ME1_C
Rg10	net037#6	net037#7	6.835e-03	$ME1_C
Rg11	net037#5	net037#6	    2.5000	$ME1_C
Rg12	avC3#9	avC3#10	   18.6250	$ME1_C
Rg13	avC3#11	avC3#12	    3.3110	$ME1_C
Rg14	avC3#12	avC3#14	    0.6277	$ME1_C
Rg15	avC3#12	avC3#11	   15.0317	$ME1_C
Rg16	avC3#14	avC3#15	    7.0310	$ME1_C
Rg17	avC3#11	avC3#12	   15.0000	$ME1_C
Rg18	avC3#13	avC3#14	   15.0000	$ME1_C
Rg19	y#1	y#2	    9.1756	$ME1_C
Rg20	net017	net017#3	   15.7775	$ME1_C
Rg21	net017#3	net017#2	   15.0214	$ME1_C
Rg22	net017#2	net017#3	   15.0000	$ME1_C
Rg23	avC3#20	avC3#21	    9.2591	$ME1_C
Rg24	avC3#23	avC3#24	   18.6257	$ME1_C
Rg25	b#12	b#9	   12.6791	$ME1_C
Rg26	net013#2	net013#3	4.126e-02	$ME1_C
Rg27	net013	net013#2	   15.0000	$ME1_C
Rg28	avC3#27	avC3#28	1.087e-02	$ME1_C
Rg29	avC3#29	avC3#30	1.097e-02	$ME1_C
Rg30	avC3#28	avC3#29	5.133e-02	$ME1_C
Rg31	avC3#32	avC3#34	1.213e-02	$ME1_C
Rg32	avC3#34	avC3#35	9.219e-03	$ME1_C
Rg33	avC3#35	avC3#36	5.774e-02	$ME1_C
Rg34	avC3#36	avC3#33	    3.2222	$ME1_C
Rg35	avC3#33	avC3#34	   15.0000	$ME1_C
Rg36	avC3#33	avC3#35	   15.0000	$ME1_C
Rg37	y#4	y#5	    9.1756	$ME1_C
Rg38	net013#5	net013#6	   15.0214	$ME1_C
Rg39	net013#6	net013#4	    0.4488	$ME1_C
Rg40	net013#5	net013#6	   15.0000	$ME1_C
Rg41	avC3#40	avC3#38	    3.1960	$ME1_C
Rg42	avC3#38	avC3#41	    3.2313	$ME1_C
Rg43	avC3#42	avC3#25	   12.3236	$ME1_C
Rg44	y	y#6	    2.3471	$ME1_C
Rg45	y#6	y#7	    1.2326	$ME1_C
Rg46	y#7	y#9	    0.4661	$ME1_C
Rg47	y#7	y#3	    0.3288	$ME1_C
Rg48	y#9	y#10	   15.9117	$ME1_C
Rg49	y#8	y#9	   15.0000	$ME1_C
Rg50	gnd#2	gnd#4	    1.6934	$ME1_C
Rg51	gnd#4	gnd#5	    0.8442	$ME1_C
Rg52	gnd#5	gnd	    0.1725	$ME1_C
Rg53	gnd	gnd#6	    1.2492	$ME1_C
Rg54	gnd#6	gnd#8	    0.3960	$ME1_C
Rg55	gnd#4	gnd#10	    0.4339	$ME1_C
Rg56	gnd#5	gnd#12	    0.3960	$ME1_C
Rg57	gnd#6	gnd#14	    1.5397	$ME1_C
Rg58	gnd#14	gnd#13	   15.0000	$ME1_C
Rg59	gnd#7	gnd#8	   15.0000	$ME1_C
Rg60	gnd#9	gnd#10	   15.0000	$ME1_C
Rg61	gnd#11	gnd#12	   15.0000	$ME1_C
Rg62	gnd#13	gnd#14	   15.0000	$ME1_C
Rg64	avC3#54	avC3#56	    1.5100	$ME1_C
Rg65	avC3#56	avC3#16	    0.4662	$ME1_C
Rg67	avC3#16	avC3#58	    0.5095	$ME1_C
Rg68	avC3#58	avC3#59	    0.2892	$ME1_C
Rg69	avC3#59	avC3#60	1.941e-03	$ME1_C
Rg70	avC3#54	avC3#62	    1.5784	$ME1_C
Rg71	avC3#62	avC3#61	   15.0000	$ME1_C
Rg72	avC3#56	avC3#6	    4.0778	$ME1_C
Rg73	avC3#16	avC3#63	    2.8558	$ME1_C
Rg74	avC3#60	avC3#22	    0.9231	$ME1_C
Rg75	avC3#22	avC3#64	    2.7591	$ME1_C
Rg76	avC3#6	avC3#66	    0.1851	$ME1_C
Rg77	avC3#66	avC3#65	   15.0000	$ME1_C
Rg78	avC3#53	avC3#54	   15.0000	$ME1_C
Rg79	avC3#53	avC3#54	   15.0000	$ME1_C
Rg80	avC3#57	avC3#58	    3.0000	$ME1_C
Rg81	avC3#57	avC3#59	   15.0000	$ME1_C
Rg82	avC3#57	avC3#60	   15.0000	$ME1_C
Rg83	avC3#61	avC3#62	   15.0000	$ME1_C
Rg84	avC3#65	avC3#66	   15.0000	$ME1_C
Rf1	gnd#1	gnd#2	   13.6853	$ME2_C
Rf2	avC3#6	avC3#4	    8.1013	$ME2_C
Rf3	net037#7	net037#3	    8.5907	$ME2_C
Rf4	avC3#16	avC3#9	    7.3101	$ME2_C
Rf5	y#3	y#2	    6.8428	$ME2_C
Rf6	avC3#20	avC3#22	    6.7729	$ME2_C
Rf7	avC3#25	avC3#26	    6.7689	$ME2_C
Rf8	avC3#26	avC3#15	    0.8758	$ME2_C
Rf9	avC3#26	avC3#24	    1.1107	$ME2_C
Rf10	net013#4	net013#3	   13.2525	$ME2_C
Rf11	avC3#36	avC3#38	   13.3854	$ME2_C
Rf12	y#5	y#6	    6.8782	$ME2_C
*
*       CAPACITOR CARDS
*
*
C1	avC3#41	avS50	2.45846e-16
C2	avC5	avC3#64	2.12843e-17
C3	avC3#9	avC9	1.19985e-17
C4	net013#3	gnd#13	3.46515e-17
C5	y#10	avC3#23	3.74297e-17
C6	net037#7	avC3	1.40129e-16
C7	avC3#41	y#4	8.20864e-18
C8	b#2	avC5	9.04944e-18
C9	net013#3	b#14	7.31375e-18
C10	y#6	avC3#40	5.55662e-17
C11	b#5	avC3#61	3.24078e-17
C12	net017	gnd#13	2.40773e-17
C13	gnd#3	avC3#47	4.36239e-17
C14	avC8	avC3#51	1.72906e-16
C15	avC3#25	gnd#13	9.26838e-17
C16	y#8	avC3#24	1.31714e-17
C17	avC3#36	avC7	1.32677e-17
C18	b#12	y#10	3.48339e-17
C19	avC3#26	gnd#13	4.12766e-17
C20	y#2	avC5	4.89256e-18
C21	y#10	gnd#13	3.50686e-17
C22	net037#4	b#10	3.0621e-17
C23	net037#8	b#12	8.60133e-18
C24	avC3#4	gnd#3	1.01054e-16
C25	b#9	gnd#13	1.55212e-16
C26	net013	b#12	3.41107e-18
C27	avC3#26	y#2	5.56163e-18
C28	net017#2	gnd#13	4.42659e-17
C29	b#2	net037#5	7.21757e-18
C30	gnd#1	b	1.33017e-16
C31	avS52	avC3#61	2.71536e-17
C32	b#3	avC5	5.81239e-18
C33	b#10	gnd#9	4.34343e-17
C34	b	gnd#13	2.03455e-16
C35	avC3#27	avC8	1.82346e-16
C36	avC3#24	gnd#13	3.22916e-17
C37	avC3#26	avC9	1.57508e-17
C38	net037#7	b#11	2.93372e-17
C39	net013#4	y#6	6.13314e-18
C40	b#7	avC3#46	1.01079e-17
C41	avC10	avC3#11	2.90707e-16
C42	avC3#52	avC9	2.50431e-16
C43	net037#8	gnd#13	4.83616e-16
C44	net037	b#10	4.32354e-17
C45	y	gnd#13	3.65988e-16
C46	net013#4	y#10	5.86776e-17
C47	net013#3	gnd#7	4.71498e-17
C48	avC3#38	y#5	1.10276e-16
C49	b#9	net037#8	1.00557e-16
C50	y#3	avC3#64	3.22121e-17
C51	avS50	net037#10	3.35692e-17
C52	avC3#31	y#6	3.8331e-17
C53	gnd#7	net013#5	2.1511e-17
C54	avC3#56	gnd#13	1.71318e-15
C55	avC3#19	gnd#13	1.68061e-16
C56	y#6	avC3#41	4.58897e-17
C57	b#9	avC3#19	9.30316e-18
C58	avC3#13	gnd#13	7.48501e-17
C59	avC3#56	avC10	1.87753e-15
C60	net037#7	b#2	2.2608e-17
C61	y#3	b#7	6.51617e-18
C62	net037#12	b#7	8.23438e-18
C63	net013#3	y#10	8.96915e-19
C64	b#5	avC3#21	2.29049e-16
C65	gnd#3	avC3#13	2.88635e-17
C66	avC3#36	avC8	9.68237e-18
C67	y#5	avC3#40	2.55286e-16
C68	avC3#53	avC7	1.15293e-16
C69	y#1	b#5	2.20988e-16
C70	avC3#24	y#6	5.83906e-17
C71	y#10	net013#5	3.7835e-17
C72	avC3#56	avC8	1.87045e-15
C73	gnd#7	net037#8	5.53348e-18
C74	net013#4	avC3#31	8.93208e-18
C75	avC5	y#3	1.86654e-17
C76	avC5	net037#5	1.07625e-17
C77	avC3#37	gnd#13	2.23562e-17
C78	avC3#42	avC8	1.78358e-16
C79	gnd#4	net037#3	1.35171e-17
C80	net037#3	b#3	3.20467e-17
C81	avS52	b#5	3.35577e-17
C82	avC3#36	avC9	3.74026e-18
C83	avC3#10	gnd#13	1.74275e-16
C84	avS52	y#1	2.21055e-16
C85	net013#4	b#13	5.14898e-17
C86	net037#8	b#7	1.62004e-17
C87	net037#8	net013	2.11718e-18
C88	net037#10	avC3#39	5.52073e-18
C89	y#10	avC3#24	5.39639e-17
C90	net013#3	b#13	1.08508e-17
C91	avC3#37	net013#5	4.96382e-17
C92	b#14	gnd#13	3.44423e-17
C93	avC3#64	avS52	2.08925e-16
C94	avC3#42	avC9	3.72873e-16
C95	avC3#25	avC7	2.86954e-17
C96	gnd#7	net013	1.20443e-18
C97	avC3#23	y#6	2.26447e-17
C98	y#10	avC3#37	4.89371e-17
C99	gnd#9	b#3	2.73581e-17
C100	avC3#24	y#5	4.18663e-17
C101	y#3	gnd#13	1.63624e-17
C102	avC8	avC3#44	4.62041e-18
C103	gnd#6	b#14	6.03793e-18
C104	avC3#41	y#5	2.57848e-16
C105	avC3#9	avC10	2.96564e-18
C106	gnd#6	net013#3	1.64672e-17
C107	avC3#46	gnd#13	1.95182e-17
C108	avC3#4	net037#7	1.48582e-17
C109	gnd#6	net013	1.299e-18
C110	avC3#57	avC9	2.22942e-16
C111	avC3#24	y#7	4.16565e-17
C112	b#14	gnd#7	5.74008e-17
C113	b#2	gnd#13	2.87157e-17
C114	avC3#9	gnd#13	4.05605e-17
C115	avC3#44	gnd#13	2.2385e-16
C116	net037#3	b#10	4.75489e-18
C117	net037#12	gnd#13	2.55696e-17
C118	b#1	net037#5	3.35494e-17
C119	net013#4	avC3#41	3.59228e-18
C120	net013	b#14	4.14747e-17
C121	avC3#56	avC9	1.87232e-15
C122	b#1	net037#7	7.65127e-17
C123	avC3#53	avC8	1.17461e-16
C124	b#3	gnd#13	1.82925e-16
C125	avC3#44	avS50	5.94763e-18
C126	net037#7	avC5	3.21684e-16
C127	net013#4	avC3#23	7.21825e-19
C128	avC3#15	gnd#13	7.34897e-17
C129	avC3#47	gnd#13	3.6631e-17
C130	y#7	avC3#20	3.29872e-17
C131	net017#2	y#3	1.727e-17
C132	net037#7	b#8	1.72596e-17
C133	avC5	b#7	3.12653e-18
C134	net013#4	b#12	3.26096e-17
C135	avC10	avC3#48	1.96257e-16
C136	avC3#61	avC8	2.44803e-17
C137	avC3#25	avC8	4.42124e-17
C138	b#8	avC3	6.22768e-17
C139	net037#7	gnd#13	1.59929e-17
C140	net013#3	b#12	3.51734e-17
C141	b#10	gnd#13	2.48051e-17
C142	avC9	avC3#44	6.94829e-18
C143	avC3#4	b#1	1.10006e-17
C144	avC9	avC3#53	1.10794e-16
C145	avC3#8	gnd#13	1.04228e-16
C146	b#11	avC5	1.88175e-16
C147	b#8	avC5	9.21826e-17
C148	net017	b#12	8.07871e-19
C149	b#13	avC3#37	8.45925e-18
C150	avC3	gnd#3	1.48062e-17
C151	net037#3	gnd#13	5.10188e-17
C152	avC3#38	net037#10	2.4289e-17
C153	gnd#1	avC3#4	6.8058e-17
C154	avC3#24	b#12	6.66359e-18
C155	avC3#39	gnd#13	9.36247e-17
C156	y#5	net037#10	3.18726e-17
C157	net037#5	b#11	1.61129e-16
C158	avC3#19	b#5	1.93414e-17
C159	avC5	avC3#13	1.06137e-17
C160	avC3#57	gnd#13	2.49903e-17
C161	avC9	avC3#61	3.21941e-17
C162	avC3#26	y#5	1.34246e-17
C163	y#2	avC3#24	1.6729e-17
C164	net013#4	b#9	1.02829e-18
C165	avC3#6	gnd#13	6.09965e-16
C166	y#6	avS50	9.74381e-18
C167	y#7	gnd#13	5.1629e-17
C168	avC3#31	gnd#13	9.63585e-17
C169	avC3#6	avC10	4.4957e-17
C170	avS52	avC3#10	3.9142e-18
C171	b#9	net013#3	1.20765e-17
C172	avC3#38	avS50	2.0753e-17
C173	b#1	gnd#13	2.13116e-16
C174	gnd#9	avC5	1.88129e-17
C175	avC3#20	y#2	2.92263e-16
C176	y#5	avS50	2.72528e-17
C177	net017#2	y#8	1.07525e-16
C178	gnd#2	net037#4	2.71628e-17
C179	avC3#4	gnd#13	1.68025e-16
C180	avC3#33	avC7	2.62513e-16
C181	b#13	gnd#13	1.07033e-16
C182	net013#3	net037#8	7.56234e-18
C183	avC3#25	avS50	1.04325e-18
C184	net013#5	avC3#31	2.23177e-17
C185	avC3#26	avS52	6.79971e-19
C186	net037#4	gnd#13	2.55238e-16
C187	avC3#20	avC9	6.36034e-18
C188	gnd#9	net037#4	8.48191e-17
C189	b#5	avC3#44	4.8389e-17
C190	b#8	net037#5	1.00895e-16
C191	avC7	avC3#39	7.89483e-16
C192	net037#4	b#3	5.24458e-18
C193	b#9	y#8	4.01453e-17
C194	y#3	avC3#24	1.2626e-17
C195	y#10	avC3#31	8.73775e-18
C196	b#11	avC3	2.75879e-17
C197	b#13	net013#5	8.48732e-18
C198	b#9	avC3#46	5.83785e-18
C199	avC3#64	y#1	5.89274e-18
C200	y#6	gnd#13	3.72636e-16
C201	gnd#4	net037#4	2.91036e-17
C202	net017	b#9	1.36768e-16
C203	gnd#4	net037#8	1.02161e-17
C204	gnd#7	b#13	2.22377e-17
C205	net037#12	b#9	1.71748e-17
C206	b#1	avC3	5.56584e-17
C207	avC3#22	y#2	1.78489e-16
C208	net037#10	avC3#61	4.28083e-17
C209	net017#2	b#9	1.04209e-18
C210	gnd#3	avC10	1.64457e-17
C211	avC3#40	y#4	8.20864e-18
C212	gnd#5	net037#8	1.67236e-17
C213	gnd#11	net017	3.46504e-17
C214	avS52	avC3#44	1.59638e-18
C215	avC3#46	y#8	4.06407e-17
C216	y#7	avC3#19	6.79454e-17
C217	y#2	avC3#21	7.92367e-18
C218	net013	b#13	5.47035e-18
C219	net037#8	net017	6.44405e-17
C220	avC3#20	y#1	8.66884e-18
C221	net017#2	avC3#46	5.206e-17
C222	net017#2	y#7	1.22157e-18
C223	avC3#20	b#5	3.29671e-17
C224	net037#10	avC3#40	2.54245e-16
C225	net037#8	net017#2	4.98665e-18
C226	avC3#38	gnd#13	5.44483e-17
C227	y#2	b#5	2.75208e-17
C228	avC3#56	avC7	1.87127e-15
C229	net013#5	y#6	2.3052e-17
C230	y#8	avC3#19	8.94173e-17
C231	gnd#11	net017#2	2.14557e-17
C232	y#4	net037#10	2.21035e-16
C233	net037#4	b#1	2.30235e-17
C234	avC3#53	gnd#13	1.34858e-16
C235	net037#7	gnd#3	1.45823e-17
C236	gnd#11	net037#8	2.00243e-16
C237	net037#12	net017	4.40491e-17
C238	avC3#20	avS52	2.23652e-18
C239	b#7	net017#2	4.07766e-17
C240	avC3#23	gnd#13	6.22365e-17
C241	avS50	avC3#61	3.80281e-17
C242	avC3#43	avC7	1.74959e-16
C243	avC3#32	avC7	2.43298e-17
C244	y#2	avS52	2.9154e-17
C245	net037#3	gnd#9	6.44768e-17
C246	net017#2	net037#12	1.86617e-18
C247	net013#4	net017	4.54115e-18
C248	avC5	avC3	5.76872e-18
C249	avC8	avC3#33	2.62282e-16
C250	avC3#15	y#2	1.14958e-17
C251	b#7	gnd#13	2.49199e-16
C252	avC3#65	avC10	1.72899e-17
C253	gnd#11	net037#12	4.11643e-17
C254	net017#2	avC3#19	4.4548e-17
C255	avC3#61	gnd#13	3.26354e-17
C256	avC3#22	avS52	2.27267e-17
C257	avC3#19	y#3	1.4979e-17
C258	b#12	gnd#13	1.25132e-16
C259	y#3	avS52	6.50018e-18
C260	net013#4	net017#2	6.66567e-18
C261	b#12	avC3#23	5.1389e-18
C262	net013#4	gnd#13	3.78938e-17
C263	avC3#40	avS50	1.59637e-18
C264	gnd#11	b#7	7.77456e-18
C265	avC3#15	avS52	1.12672e-18
C266	net013#3	net017	6.85144e-18
C267	net013#5	gnd#13	7.07798e-17
C268	avS50	y#4	2.21168e-16
C269	y#2	avC3#64	2.2111e-16
C270	y#5	avC3#61	6.09516e-18
C271	net013#4	avC3#37	6.83045e-18
C272	avC8	avC3#32	1.03673e-16
C273	avC3#42	gnd#13	8.96003e-17
C274	y#8	gnd#13	2.81126e-17
C275	avC3#15	b#6	2.50887e-17
C276	net017#2	b#6	2.45901e-18
C277	gnd#3	avC3#7	1.94081e-17
C278	y#2	b#6	5.32243e-18
C279	net017#2	net037#11	8.11448e-18
C280	avC5	b#6	3.4721e-17
C281	b#6	avS52	4.86504e-17
C282	avC9	avC3#16	8.22152e-17
C283	net037#11	avC3#41	1.35247e-16
C284	avC3#16	gnd#13	6.16445e-17
C285	net013#4	net037#11	1.06893e-17
C286	avC3#26	net037#11	8.70732e-18
C287	b#6	avC3#19	7.23916e-17
C288	b#6	gnd#13	3.12924e-16
C289	net037#11	avC3#23	5.08045e-17
C290	y#8	net037#11	6.49328e-17
C291	b#6	y#1	6.47821e-18
C292	avC3#24	net037#11	4.12936e-17
C293	net037#11	avC3#61	1.35693e-16
C294	y#7	net037#11	6.82396e-17
C295	avC3#31	net037#11	4.19277e-17
C296	net037#11	y#4	6.47821e-18
C297	avC3#22	b#6	2.17874e-17
C298	avC3#7	avC10	2.47754e-16
C299	net037#11	y#10	8.37364e-18
C300	avC3#19	net037#11	8.76541e-17
C301	y#3	b#6	5.22157e-17
C302	net037#11	gnd#13	4.43132e-16
C303	avC3#7	gnd#13	4.60419e-16
C304	y#7	b#6	3.64348e-17
C305	b#6	avC3#61	7.73052e-17
C306	b#6	avC3#64	1.3327e-16
C307	y#6	net037#11	9.18989e-17
C308	avC3#20	net037#11	1.33373e-17
C309	net037#11	avS50	4.86096e-17
C310	net013#5	net037#11	3.79038e-18
C311	b#9	net037#11	5.80187e-18
C312	y#5	net037#11	1.17987e-17
C313	avC3#44	net037#11	3.94804e-17
C314	gnd#2	b#1	3.13364e-18
C315	gnd#4	b#10	3.1585e-18
C316	gnd#2	b	3.95334e-18
C317	y#7	b#9	1.28091e-18
C318	y#6	b#13	2.3062e-18
C319	b#13	y#10	2.91492e-18
C320	y#7	b#5	3.55917e-18
C321	avC3#15	gnd#3	4.28091e-18
C322	gnd#1	avC3	5.40196e-18
C323	gnd#3	avC3#8	9.64537e-18
C324	net037#7	b#7	1.4217e-18
C325	net037#8	b#3	1.73951e-18
C326	net037#7	b#3	2.22014e-18
C327	net037	b#8	2.33667e-18
C328	net037#8	b#14	3.03609e-18
C329	net037#3	b#8	4.59937e-18
C330	net037#7	b#6	4.69952e-18
C331	avC3#41	b#5	1.31516e-18
C332	avC3#22	b#5	1.36637e-18
C333	b#13	avC3#31	1.86766e-18
C334	avC3#13	b#6	2.23942e-18
C335	avC3#15	b#5	2.36258e-18
C336	avC3#47	b#6	2.40339e-18
C337	avC3#4	b#11	2.53431e-18
C338	b#2	avC3	2.91954e-18
C339	b#11	avC3#47	3.06431e-18
C340	b#6	avC3#10	4.05895e-18
C341	y#3	net037#11	4.17046e-18
C342	avC8	avC3#43	1.86396e-18
C343	y#5	avC3#20	1.5187e-18
C344	y#3	avC3#20	1.73414e-18
C345	y#1	avC3#44	2.24847e-18
C346	y#4	avC3#39	2.28567e-18
C347	y#2	avC3#41	2.39233e-18
C348	y#3	avC3#61	2.62749e-18
C349	y#7	avC3#21	2.67999e-18
C350	y#2	avC3#44	3.03514e-18
C351	avC3#22	y#1	3.84853e-18
C352	y#2	avC3#19	4.07656e-18
C353	y#6	avC3#61	4.37005e-18
C354	avC3#20	avS50	5.69132e-19
C355	avC3#41	net037#10	2.41369e-18
C356	avC3#25	net037#11	2.95087e-18
C357	net037#11	avC3#37	2.97208e-18
C358	avC3#46	net037#11	4.11461e-18
C359	avC3#38	net037#11	4.65299e-18
C360	avC3#9	avS52	5.58639e-19
C361	net013#4	net037#8	5.28091e-19
C362	net037#10	gnd	7.48417e-18
C363	avS50	gnd	4.45406e-19
C364	avC3#51	gnd	3.46186e-18
C365	avC3#52	gnd	1.1357e-18
C366	b#5	gnd	3.85602e-18
C367	avS52	gnd	8.78159e-19
C368	avC3#17	gnd	1.36716e-18
C369	b#11	gnd	1.02564e-18
C370	avC3#46	gnd	1.36484e-18
C371	avC3#39	gnd	1.03802e-18
C372	avC3#31	gnd	2.67005e-19
C373	b#13	gnd	1.27809e-18
C374	avC3#32	gnd	2.84038e-19
C375	avC3#30	gnd	2.33733e-19
C376	avC3#23	gnd	1.63018e-18
C377	b#12	gnd	8.81957e-19
C378	b#9	gnd	8.98345e-18
C379	net037#8	gnd	3.18908e-17
C380	avC3#19	gnd	9.90055e-19
C381	b#2	gnd	1.44959e-18
C382	avC3#7	gnd	3.84338e-20
C383	avC3#8	gnd	1.26182e-18
C384	b#1	gnd	2.239e-18
C385	net037#4	gnd	1.07495e-18
C386	y#6	gnd	4.15616e-18
C387	avC3#38	gnd	9.0123e-18
C388	y#5	gnd	5.67906e-19
C389	net013#3	gnd	3.07999e-19
C390	avC3#25	gnd	1.64729e-18
C391	avC3#24	gnd	9.75643e-19
C392	y#2	gnd	1.35353e-18
C393	avC3#22	gnd	4.10728e-18
C394	y#3	gnd	1.59742e-18
C395	avC3#9	gnd	8.34843e-19
C396	net013#5	gnd	4.34671e-19
C397	avC7	gnd	2.60838e-18
C398	y#4	gnd	1.45291e-18
C399	avC8	gnd	5.69616e-18
C400	avC9	gnd	6.57412e-18
C401	avC3#21	gnd	1.10438e-18
C402	avC3#57	gnd	4.61037e-19
C403	avC3#64	gnd	1.16452e-18
C404	avC3#11	gnd	3.18241e-18
C405	avC5	gnd	8.2411e-18
C406	avC10	gnd	1.26182e-18
C407	net037#5	gnd	1.55146e-20
C408	y#8	gnd	4.06707e-18
C409	net017	gnd	8.75044e-18
C410	net017#2	gnd	8.07277e-18
C411	net037	gnd	7.33455e-19
C412	b#6	gnd	1.96841e-18
C413	b#7	gnd	1.39669e-18
C414	b#8	gnd	1.07495e-18
C415	avC3#26	gnd	1.99611e-18
C416	net037#11	gnd	3.36049e-18
C417	avC3#44	gnd	6.30272e-19
C418	y#7	gnd	2.80738e-19
*
*
.ENDS XNOR2X1
*
